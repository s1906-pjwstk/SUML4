���	     �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�	estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �_sklearn_version��1.3.2�ub�n_estimators�Kd�estimator_params�(hhhhhhhhhht��base_estimator��
deprecated��	bootstrap���	oob_score���n_jobs�NhK*�verbose�K �
warm_start��hN�max_samples�NhhhNhKhKhG        h�sqrt�hNhG        hG        �feature_names_in_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h+�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�Pclass��Sex��Age��SibSp��Parch��Fare��Embarked�et�b�n_features_in_�K�
n_outputs_�K�classes_�h*h-K ��h/��R�(KK��h4�i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�K�
estimator_�h	�estimators_�]�(h)��}�(hhhhhNhKhKhG        hh&hNhJf��_hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h4�f8�����R�(KhMNNNJ����J����K t�b�C              �?�t�bhQh(�scalar���hLC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hK�
node_count�M?�nodes�h*h-K ��h/��R�(KM?��h4�V64�����R�(Kh8N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples��missing_go_to_left�t�}�(h}hLK ��h~hLK��hhLK��h�h]K��h�h]K ��h�hLK(��h�h]K0��h�h4�u1�����R�(Kh8NNNJ����J����K t�bK8��uK@KKt�b�B�O                            �?z����?�           @�@              	                   �0@�x�c���?T           Ȁ@                                @�&@     ��?	             0@       ������������������������       �                     $@                                  �,@r�q��?             @                                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        
       e                    �?HT,��l�?K           H�@                                   �8@z91$UO�?X            �a@                                 s�@$��m��?             :@                                   �?r�q��?             @        ������������������������       �                      @                                �{@      �?             @        ������������������������       �                     �?                                  �4@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                  �7@z�G�z�?             4@                                 @,@�	j*D�?	             *@                                  �#@      �?              @                                  �5@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                                   �?���Q��?             @                                 �1@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        !       `                    �?�c����?H            @]@       "       S                 @�6M@4uj�w��?E            @\@       #       0                     @�DC��,�?7            �V@        $       /                    �?     ��?             0@       %       (                    �?�q�q�?             (@        &       '                   �4@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        )       *                 ���,@      �?              @        ������������������������       �                      @        +       ,                 0C�?@�q�q�?             @        ������������������������       �                      @        -       .                   �B@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        1       <                  ��@DE��2{�?,            �R@        2       5                    �?�t����?             A@        3       4                 �Y�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        6       ;                   @<@��a�n`�?             ?@       7       :                    �?ȵHPS!�?             :@       8       9                 ���@�S����?	             3@        ������������������������       �                     $@        ������������������������       ��q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        =       H                 �̌@������?            �D@        >       ?                    �?�G��l��?             5@        ������������������������       �                      @        @       G                    �?8�Z$���?	             *@       A       D                   �<@r�q��?             (@       B       C                 ��(@�����H�?             "@       ������������������������       �      �?              @        ������������������������       �                     �?        E       F                   �H@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        I       N                    �?ףp=
�?             4@       J       M                    ;@�8��8��?             (@        K       L                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        O       R                    �?      �?              @        P       Q                 03�'@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        T       _                    �?"pc�
�?             6@       U       V                    �?��s����?             5@       ������������������������       �                     *@        W       Z                    �?      �?              @        X       Y                 p�w@      �?             @       ������������������������       �                      @        ������������������������       �                      @        [       \                    C@      �?             @        ������������������������       �                     �?        ]       ^                   �H@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        a       b                    �?      �?             @        ������������������������       �                     �?        c       d                  �v6@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        f       �                    �?�V���?�            �w@        g       �                   �<@�X����?;             V@       h       y                   �8@~|z����?             �J@       i       x                 pF�'@X�Cc�?             <@       j       w                    �?      �?             0@       k       v                   �6@      �?	             (@       l       s                   �4@�eP*L��?             &@        m       r                    3@���Q��?             @       n       o                 P��@      �?             @        ������������������������       �                     �?        p       q                 ��!@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        t       u                 جJ"@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        z                        03�$@���Q��?             9@        {       |                   �9@ףp=
�?             $@        ������������������������       �                     @        }       ~                    ;@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �̌2@���Q��?             .@       �       �                     @�����H�?             "@        ������������������������       �                     @        �       �                    ;@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ��TS@r�q��?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    @@�#-���?            �A@        �       �                     @z�G�z�?             $@        ������������������������       �                     @        �       �                 @3#%@      �?             @        ������������������������       �                     �?        �       �                 ��y.@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?`2U0*��?             9@       ������������������������       �                     ,@        �       �                     @�C��2(�?	             &@       ������������������������       �                     "@        �       �                    D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ��$:@<�f~�?�             r@       �       �                 ��@\�$����?�             m@        �       �                 ��@��<b�ƥ?             G@        �       �                 ��@P���Q�?             4@       ������������������������       �                     3@        ������������������������       �                     �?        ������������������������       �                     :@        �       �                   �<@h�O,��?w            `g@       �       �                 �1@@4և���?D            �X@        �       �                   �9@      �?              @       ������������������������       �                     @        ������������������������       �                     @        �       �                   �4@`Ӹ����??            �V@        �       �                 pf� @      �?	             (@       �       �                   �3@      �?             @        ������������������������       �      �?              @        �       �                 P�@      �?             @        ������������������������       �                     �?        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   �;@�(�Tw�?6            �S@        �       �                   �:@������?             B@       ������������������������       �                    �A@        ������������������������       �                     �?        ������������������������       �                     E@        �       �                 @3�@4\�����?3            @V@        �       �                 �?�@�	j*D�?             :@        �       �                   �?@$�q-�?             *@        ������������������������       �                     "@        �       �                   �A@      �?             @       �       �                   �@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   @A@��
ц��?             *@        ������������������������       �                     @        �       �                    �?���Q��?             $@       �       �                   �D@և���X�?             @       ������������������������       ����Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   @@@�����?(            �O@        �       �                   �7@������?             .@       �       �                   �=@d}h���?
             ,@        �       �                     @�q�q�?             @        ������������������������       �                     @        �       �                 ���"@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ��i @      �?              @        �       �                    ?@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    M@ �q�q�?             H@       �       �                     @��<b�ƥ?             G@       �       �                   �*@XB���?             =@        �       �                 `fF)@      �?	             0@        ������������������������       �                     @        �       �                   �F@$�q-�?             *@       �       �                   @D@؇���X�?             @        ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �        	             *@        ������������������������       �        	             1@        �       �                   �P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�q�q�?#            �L@       �       �                     @�K��&�?            �E@       �       �                     �?b�2�tk�?             B@       �       �                   @>@4���C�?            �@@       �       �                 03k:@�ՙ/�?             5@        ������������������������       �                      @        �       �                   �Q@D�n�3�?             3@       �       �                 `f�;@      �?             0@       �       �                   �K@��
ц��?             *@       �       �                   @G@�<ݚ�?             "@       �       �                   @B@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   �<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    @@�8��8��?             (@        �       �                   �J@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    ;@և���X�?             @        ������������������������       �                      @        �       �                    >@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �                           �?@4և���?             ,@       �                        03�U@�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        ������������������������       �                      @              >                   @s8?U��?o            �e@                             �Q��?k�q��?m            @e@        ������������������������       �                     @                                  @�W����?j            �d@                                �?N�zv�?6             V@                                @XB���?"             M@        	      
                ��1V@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      K@                                  @�������?             >@                                �?R�}e�.�?             :@                             �̾w@���N8�?             5@                                �?�S����?             3@        ������������������������       �                     $@                                 �?�q�q�?             "@        ������������������������       �                     �?                                 :@      �?              @        ������������������������       �                     �?                                 D@؇���X�?             @                               x�C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @                                 -@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @               5                `v�6@|�i���?4             S@       !      &                  �*@X��ʑ��?            �E@        "      %                   <@      �?             (@       #      $                   �?ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                      @        '      4                    @�P�*�?             ?@       (      -                   �?П[;U��?             =@        )      ,                   3@�q�q�?             @        *      +                   #@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        .      /                `ff.@�û��|�?             7@        ������������������������       �                     @        0      1                   �?      �?             2@        ������������������������       �                     @        2      3                   #@      �?             (@        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                      @        6      7                   �?Pa�	�?            �@@        ������������������������       �        
             .@        8      9                   �?�X�<ݺ?             2@        ������������������������       �                      @        :      =                   @      �?             0@        ;      <                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ,@        ������������������������       �                     @        �t�b�values�h*h-K ��h/��R�(KM?KK��h]�B�       �{@     �p@     �v@     �e@      @      &@              $@      @      �?      �?      �?              �?      �?              @             pv@     @d@     �T@     �N@      "@      1@      @      �?       @              @      �?      �?               @      �?              �?       @              @      0@      @      "@      �?      @      �?      @      �?                      @              @      @       @      �?       @      �?                       @       @                      @     @R@      F@      R@     �D@      Q@      7@      "@      @      @      @      �?      @              @      �?              @      @               @      @       @       @               @       @               @       @              @             �M@      0@      >@      @       @      �?              �?       @              <@      @      7@      @      0@      @      $@              @      @      @              @              =@      (@      &@      $@               @      &@       @      $@       @       @      �?      @      �?      �?               @      �?              �?       @              �?              2@       @      &@      �?      �?      �?              �?      �?              $@              @      �?      �?      �?      �?                      �?      @              @      2@      @      1@              *@      @      @       @       @       @                       @       @       @      �?              �?       @               @      �?                      �?      �?      @              �?      �?       @      �?                       @     Pq@     @Y@      <@      N@      9@      <@      $@      2@      $@      @      @      @      @      @      @       @       @       @              �?       @      �?       @                      �?      �?               @      @              @       @              �?              @                      (@      .@      $@      "@      �?      @              @      �?              �?      @              @      "@      �?       @              @      �?      @      �?                      @      @      �?      @                      �?      @      @@       @       @              @       @       @      �?              �?       @               @      �?              �?      8@              ,@      �?      $@              "@      �?      �?              �?      �?              o@     �D@     `j@      6@     �F@      �?      3@      �?      3@                      �?      :@             �d@      5@     �V@      @      @      @      @                      @     �U@      @      "@      @      @      @      �?      �?       @       @      �?              �?       @      �?                       @      @             @S@      �?     �A@      �?     �A@                      �?      E@             �R@      ,@      2@       @      (@      �?      "@              @      �?      �?      �?              �?      �?               @              @      @              @      @      @      @      @      @       @               @      @             �L@      @      &@      @      &@      @      @       @      @              �?       @      �?                       @      @      �?       @      �?       @                      �?      @                      �?      G@       @     �F@      �?      <@      �?      .@      �?      @              (@      �?      @      �?      @               @      �?      @              *@              1@              �?      �?              �?      �?              C@      3@      9@      2@      6@      ,@      3@      ,@       @      *@               @       @      &@       @       @      @      @       @      @       @       @      �?       @      �?                      @      @               @      �?              �?       @                      @      &@      �?      @      �?              �?      @               @              @              @      @               @      @       @      @                       @      *@      �?      &@      �?      &@                      �?       @             �T@      W@     �S@      W@              @     �S@     �U@      9@     �O@       @      L@       @       @               @       @                      K@      7@      @      3@      @      0@      @      0@      @      $@              @      @              �?      @       @              �?      @      �?      �?      �?      �?                      �?      @                       @      @       @               @      @              @             �J@      7@      5@      6@      @      "@      �?      "@      �?                      "@       @              2@      *@      0@      *@       @      @       @      �?              �?       @                      @      ,@      "@      @              "@      "@              @      "@      @              @      "@               @              @@      �?      .@              1@      �?       @              .@      �?      �?      �?      �?                      �?      ,@              @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�=�KhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B@C         V                    �?��!h
��?�           @�@               O                 p�H@�Ee@���?�            �n@              H                    @�F ���?r            �d@                                  !@��Sݭg�?l            �c@        ������������������������       �                     3@                                    @�5Q^�u�?`             a@               
                     �?���N8�?!             E@               	                   �H@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                  @4@ ���J��?            �C@        ������������������������       �                     4@                                  �;@�}�+r��?             3@                                  �7@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        	             $@               '                    �?���Q��??            �W@                                  �6@��R[s�?            �A@                                 s�@����X�?             @                                03�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @               "                    �?؇���X�?             <@              !                    �?�8��8��?             8@                                pF @�r����?
             .@                               ���@@4և���?	             ,@        ������������������������       �                     @                                �&B@ףp=
�?             $@       ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@        #       &                 `�@1@      �?             @       $       %                   �<@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        (       G                 ���4@�������?'             N@       )       F                    C@Fx$(�?             I@       *       ;                 `f�%@�I� �?             G@       +       :                    �?X�<ݚ�?             ;@       ,       3                 pf� @
j*D>�?             :@       -       .                 ���@      �?             0@        ������������������������       �                     @        /       2                   �9@�	j*D�?             *@       0       1                   �6@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        4       7                  �#@�z�G��?             $@       5       6                   �;@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        8       9                 �[$@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        <       =                    �?�S����?             3@        ������������������������       �                     @        >       C                    �?�θ�?	             *@       ?       @                 @3�/@z�G�z�?             $@        ������������������������       �                     @        A       B                    ;@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        D       E                 03S1@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     $@        I       J                 ���3@"pc�
�?             &@        ������������������������       �                     �?        K       N                    @ףp=
�?             $@        L       M                    @      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        P       U                     @�kb97�?3            @S@       Q       R                    �?��
���?1            �R@       ������������������������       �        *            �O@        S       T                     @r�q��?             (@        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �                      @        W       ^                    $@tk~X��?           @}@        X       Y                    �?�X����?             6@        ������������������������       �                      @        Z       [                    @      �?             4@       ������������������������       �        	             ,@        \       ]                    @r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        _       �                 ���<@P�@�I�?           �{@       `       {                    �?�O�5Ҫ�?�            `v@        a       z                 ��d5@�GN�z�?             F@       b       y                    �?�E��ӭ�?             B@       c       d                     @�t����?             A@        ������������������������       �                      @        e       p                    ;@      �?             @@        f       g                 ��y@      �?             (@        ������������������������       �                      @        h       i                    /@���Q��?             $@        ������������������������       �                     �?        j       k                 ���@�q�q�?             "@        ������������������������       �                     @        l       o                 xF*@      �?             @       m       n                    5@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        q       x                   �=@ףp=
�?             4@       r       s                 ���@8�Z$���?
             *@        ������������������������       �                     @        t       u                   @@      �?              @       ������������������������       �z�G�z�?             @        v       w                   �<@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        |       �                    �?�Z��=��?�            �s@       }       �                     @p�"�0�?�            �r@        ~       �                   @N@h��@D��?3            �Q@              �                    �?t�e�í�?1            �P@        ������������������������       �                      @        �       �                   �@@$�q-�?0            @P@       �       �                    &@��?^�k�?            �A@        �       �                     �?�C��2(�?	             &@        ������������������������       �                     �?        �       �                    @ףp=
�?             $@        ������������������������       �                     @        �       �                   �1@؇���X�?             @        ������������������������       �                      @        �       �                   �6@z�G�z�?             @        ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     8@        �       �                 ��$:@�r����?             >@       �       �                    �?HP�s��?             9@       �       �                   �*@ףp=
�?             4@       �       �                   �F@8�Z$���?
             *@       �       �                    @�<ݚ�?             "@        ������������������������       �                      @        �       �                   @D@����X�?             @       �       �                   @B@z�G�z�?             @       ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �E@���Q��?             @        ������������������������       �                     �?        �       �                    H@      �?             @        ������������������������       �                      @        �       �                   �J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �P@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �:@l=fՆ�?�            `l@        �       �                   �5@xdQ�m��?0            @T@       �       �                    �?�*/�8V�?            �G@       �       �                 ��Y @�q��/��?             G@       �       �                 �?$@�חF�P�?             ?@        ������������������������       �                     ,@        �       �                 �1@�t����?             1@        ������������������������       �                      @        �       �                 @3�@z�G�z�?
             .@        ������������������������       �                      @        �       �                   �3@և���X�?             @       �       �                   �1@���Q��?             @        ������������������������       �      �?              @        ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     .@        ������������������������       �                     �?        ������������������������       �                     A@        �       �                    �?b<g���?S            @b@       �       �                  s�@:	��ʵ�?L            �`@        �       �                 P�@г�wY;�?             A@        �       �                   �;@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     8@        �       �                    �?�9�z���?:            @Y@        �       �                   �=@�J�4�?             9@       �       �                 ��(@z�G�z�?
             4@       ������������������������       ��	j*D�?             *@        ������������������������       �                     @        ������������������������       �                     @        �       �                   �;@      �?-             S@        ������������������������       �                     @        �       �                   �@��oh���?,            @R@        �       �                 ��L@��
ц��?             *@       �       �                   �=@���|���?             &@       �       �                 �?$@�q�q�?             @       ������������������������       �z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                 �?�@r�q��?&             N@        ������������������������       �                     3@        �       �                 @3�@���?            �D@        ������������������������       �                     @        �       �                   @@@4?,R��?             B@       �       �                    ?@�GN�z�?             6@       �       �                 ��) @��s����?             5@       ������������������������       �                     *@        �       �                   �<@      �?              @       �       �                 �̜!@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                 ���"@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        	             ,@        ������������������������       �                     &@        ������������������������       �        
             0@        �       �                   �8@�X���?4             V@        ������������������������       �                     $@        �       �                    �?�n_Y�K�?-            �S@        �       �                   �G@� �	��?             9@       �       �                    �?�G�z��?             4@       �       �                 ���=@��.k���?
             1@        ������������������������       �                     @        �       �                    �?և���X�?	             ,@       �       �                    �?      �?             @       �       �                   �;@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   �:@      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �;@�q����?            �J@        ������������������������       �                     @        �                           �? \� ���?            �H@       �                          �?�E��ӭ�?             B@       �       �                    @@r٣����?            �@@        ������������������������       �                     @        �       �                 ��4U@\-��p�?             =@       �       �                    �?`2U0*��?             9@       ������������������������       �                     3@        �       �                  x�N@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �                          �B@      �?             @        ������������������������       �                      @                                 �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                 �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                              p�O@8�Z$���?	             *@             	                0��G@�q�q�?             @        ������������������������       �                     @        
                         >@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �t�bh�h*h-K ��h/��R�(KMKK��h]�B�       �z@     �q@     �J@     �g@     �H@     �]@      D@      ]@              3@      D@     @X@       @      D@      �?       @               @      �?              �?      C@              4@      �?      2@      �?       @      �?                       @              $@      C@     �L@      "@      :@      @       @      �?       @      �?                       @      @              @      8@       @      6@       @      *@      �?      *@              @      �?      "@      �?      @               @      �?                      "@       @       @       @      �?       @                      �?              �?      =@      ?@      3@      ?@      .@      ?@      (@      .@      &@      .@      @      (@              @      @      "@      @      @              @      @                      @      @      @      @      �?      @                      �?      �?       @               @      �?              �?              @      0@              @      @      $@       @       @              @       @      @       @                      @      �?       @      �?                       @      @              $@              "@       @              �?      "@      �?      @      �?      @                      �?      @              @     @R@       @     @R@             �O@       @      $@       @                      $@       @             �w@     �V@      @      .@       @              @      .@              ,@      @      �?      @                      �?      w@      S@     �s@      G@      A@      $@      :@      $@      8@      $@               @      8@       @      @      @       @              @      @      �?              @      @              @      @      @      @       @               @      @                      �?      2@       @      &@       @      @              @       @      @      �?       @      �?       @                      �?      @               @               @             `q@      B@     `p@      B@      P@      @      O@      @       @              N@      @      A@      �?      $@      �?      �?              "@      �?      @              @      �?       @              @      �?       @      �?       @              8@              :@      @      7@       @      2@       @      &@       @      @       @       @              @       @      @      �?       @      �?       @              �?      �?      @              @              @              @       @              �?      @      �?       @              �?      �?              �?      �?               @       @               @       @             �h@      =@      S@      @      E@      @     �D@      @      :@      @      ,@              (@      @               @      (@      @       @              @      @       @      @      �?      �?      �?       @       @              .@              �?              A@             �^@      8@     �[@      8@     �@@      �?      "@      �?              �?      "@              8@             �S@      7@      5@      @      0@      @      "@      @      @              @             �L@      3@              @     �L@      0@      @      @      @      @       @      @      �?      @      �?              @                       @      I@      $@      3@              ?@      $@              @      ?@      @      1@      @      1@      @      *@              @      @       @       @               @       @               @       @       @                       @              �?      ,@              &@              0@              M@      >@      $@              H@      >@      &@      ,@      &@      "@       @      "@              @       @      @      @      @      @      �?              �?      @                       @      @      @              @      @              @                      @     �B@      0@              @     �B@      (@      :@      $@      9@       @              @      9@      @      8@      �?      3@              @      �?              �?      @              �?      @               @      �?      �?              �?      �?              �?       @      �?                       @      &@       @      @       @      @              �?       @      �?                       @      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ\bshG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM%huh*h-K ��h/��R�(KM%��h|�B@I                             �?z��Y�)�?�           @�@                                   @$�q-�?             *@       ������������������������       �                     (@        ������������������������       �                     �?                               ��gS@HC[X;��?�           ؅@                                 @��|��?�           X�@              ^                    �?v�����?p           �@               Q                    �?���!pc�?t            `g@       	                            @x��}�?b            �d@        
                           �?0��P�?0            �T@                               03[=@85�}C�?&            �N@                               ���;@���H��?             E@                                  �?������?            �D@                               ��Y)@`Jj��?             ?@        ������������������������       �                     *@                                   :@�����H�?             2@                                  �5@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     ,@                                  �6@z�G�z�?             $@                                   �?���Q��?             @        ������������������������       �                     �?                                  �<@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     3@        ������������������������       �        
             5@               0                 pF @|jq��?2            �T@                '                    �?��� ��?             ?@        !       "                    �?      �?
             0@        ������������������������       �                     @        #       &                    4@�C��2(�?             &@        $       %                    1@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        (       )                    0@z�G�z�?             .@        ������������������������       �                     �?        *       /                   �;@؇���X�?
             ,@       +       ,                 P�@$�q-�?	             *@       ������������������������       �                     @        -       .                   �8@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        1       6                    �?
j*D>�?             J@        2       3                    �?�<ݚ�?             "@        ������������������������       �                     @        4       5                    �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        7       L                   �@@v ��?            �E@       8       K                    @b�2�tk�?             B@       9       J                    �?j���� �?             A@       :       ;                    �?����e��?            �@@        ������������������������       �                     @        <       A                    3@����X�?             <@        =       @                   �&@r�q��?             @       >       ?                   �#@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        B       C                 ��&@��2(&�?             6@        ������������������������       �                      @        D       I                   �>@d}h���?             ,@       E       H                    �?�q�q�?             "@       F       G                    ;@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        M       P                   `1@؇���X�?             @       N       O                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        R       W                   �5@�eP*L��?             6@        S       V                    �?���!pc�?             &@        T       U                    !@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        X       Y                     @���|���?
             &@        ������������������������       �                     @        Z       ]                    �?z�G�z�?             @       [       \                    :@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        _       �                    �?�t����?�            px@       `       �                 �?�@�C���?�            �u@        a       v                   �9@�d���Ҹ?\             a@        b       u                 �1@      �?             D@       c       t                    �?r�q��?             >@       d       i                    �?�+$�jP�?             ;@        e       f                 ���@z�G�z�?             @        ������������������������       �                     @        g       h                    5@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        j       q                 �?$@"pc�
�?             6@       k       l                    7@�����H�?             2@       ������������������������       �        	             &@        m       n                   �8@����X�?             @        ������������������������       �                     �?        o       p                 @33@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        r       s                   �6@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     $@        w       ~                    �?`�E���?>            @X@        x       }                   �>@���7�?             6@       y       z                 ���@@4և���?
             ,@        ������������������������       �                     @        {       |                   @@�����H�?             "@       ������������������������       �z�G�z�?             @        ������������������������       �                     @        ������������������������       �                      @               �                     @�}��L�?/            �R@        ������������������������       �                     &@        �       �                    �?     ��?(             P@        ������������������������       �                     4@        �       �                    =@`���i��?             F@       �       �                    ;@`2U0*��?             9@        ������������������������       �                     @        �       �                  sW@�}�+r��?             3@        �       �                 pf�@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     3@        �       �                    �?�r�.kx�?�            @j@        �       �                    �?�q�q�?             8@       �       �                     �?�z�G��?             4@        �       �                 ���<@�q�q�?             @        ������������������������       �                     @        �       �                 `f�B@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                     @����X�?	             ,@        �       �                 ���,@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �*@�z�G��?             $@        ������������������������       �                     �?        �       �                   �2@�<ݚ�?             "@        ������������������������       �                     @        �       �                    �?���Q��?             @       �       �                    ;@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �>@X��Oԣ�?v            @g@       �       �                 @3�@,Z0R�?G             ]@        ������������������������       �                     �?        �       �                    &@���^���?F            �\@       �       �                    �?\#r��?&            �N@       �       �                   �0@ףp=
�?%             N@        �       �                 �̌"@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                     @��ϭ�*�?#             M@        �       �                   �5@r�q��?             (@        ������������������������       ����Q��?             @        ������������������������       �                     @        �       �                   �:@���.�6�?             G@        ������������������������       �                     8@        �       �                 pf� @��2(&�?             6@       ������������������������       �                     *@        �       �                   �;@�q�q�?             "@        ������������������������       �                      @        �       �                   �<@؇���X�?             @       ������������������������       �                     @        �       �                 ���"@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    :@ 7���B�?              K@        ������������������������       �                     >@        �       �                   �;@�8��8��?             8@        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   @<@P���Q�?             4@       �       �                   �+@      �?
             0@        ������������������������       �                     �?        ������������������������       �        	             .@        ������������������������       �                     @        �       �                 @3�@b�h�d.�?/            �Q@        �       �                   �?@�q�q�?             @        ������������������������       �                      @        �       �                   �D@      �?             @       �       �                   �A@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ��$:@      �?*             P@       �       �                     @�}�+r��?             C@       �       �                   �E@$�q-�?             :@        �       �                   @D@8�Z$���?	             *@       �       �                    1@�C��2(�?             &@       �       �                   �'@؇���X�?             @        ������������������������       �                      @        ������������������������       �z�G�z�?             @        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �        	             *@        ������������������������       �                     (@        �       �                   �J@�θ�?             :@       �       �                   �G@�q�q�?             2@       �       �                   �E@�8��8��?             (@        �       �                    �?z�G�z�?             @        �       �                 �!2C@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                     �?�GN�z�?             F@        ������������������������       �                     @        �       �                   �3@��Sݭg�?            �C@        �       �                     @     ��?             0@        ������������������������       �                      @        �       �                 �=.@      �?
             ,@       �       �                    �?����X�?             @        �       �                   @7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 P��)@      �?             @       �       �                    &@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?����X�?             @        ������������������������       �                      @        ������������������������       �                     @        �                            @�nkK�?             7@       �       �                    �?�C��2(�?             &@       �       �                    &@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     (@                                 �?��Y��]�?            �D@                              pf�C@�IєX�?             1@                              ��T?@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     8@        	                         �?     ��?.             T@        
                         �?�?�'�@�?             C@                                =@�t����?             1@                              `��Z@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                     5@                                 �?�G��l��?             E@                                �?`�Q��?             9@        ������������������������       �                     .@                              ��Q^@z�G�z�?	             $@                             Ј�U@�����H�?             "@        ������������������������       �                     @                                 �?      �?             @                               �@@�q�q�?             @        ������������������������       �                     �?                              @�pX@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?                                  �?�t����?             1@        ������������������������       �                     $@        !      "                   �?����X�?             @        ������������������������       �                     @        #      $                   5@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �t�b��-     h�h*h-K ��h/��R�(KM%KK��h]�BP       �|@     @o@      �?      (@              (@      �?             �|@     �m@     @{@     �f@     �x@     �f@     �I@      a@     �C@     �_@      @     @S@      @      L@      @     �B@      @     �B@       @      =@              *@       @      0@       @       @               @       @                      ,@       @       @       @      @              �?       @       @       @                       @              @      �?                      3@              5@      A@     �H@      @      ;@      �?      .@              @      �?      $@      �?      @              @      �?                      @      @      (@      �?               @      (@      �?      (@              @      �?      @      �?                      @      �?              >@      6@      @       @      @              @       @      @                       @      7@      4@      6@      ,@      4@      ,@      4@      *@              @      4@       @      �?      @      �?       @               @      �?                      @      3@      @       @              &@      @      @      @      @      @      @                      @      @              @                      �?       @              �?      @      �?       @               @      �?                      @      (@      $@       @      @      �?      @              @      �?              @              @      @              @      @      �?       @      �?              �?       @               @             �u@      G@     ps@      B@     @`@      @     �A@      @      9@      @      6@      @      @      �?      @              �?      �?              �?      �?              2@      @      0@       @      &@              @       @              �?      @      �?              �?      @               @       @               @       @              @              $@             �W@       @      5@      �?      *@      �?      @               @      �?      @      �?      @               @             �R@      �?      &@             �O@      �?      4@             �E@      �?      8@      �?      @              2@      �?      @      �?      @                      �?      &@              3@             �f@      =@      0@       @      ,@      @      @       @      @              �?       @               @      �?              $@      @      @      �?              �?      @              @      @              �?      @       @      @              @       @       @       @               @       @              �?               @       @       @                       @     �d@      5@     �Z@      "@              �?     �Z@       @     �K@      @      K@      @      �?      �?              �?      �?             �J@      @      $@       @      @       @      @             �E@      @      8@              3@      @      *@              @      @               @      @      �?      @               @      �?       @                      �?      �?              J@       @      >@              6@       @      @      �?      @                      �?      3@      �?      .@      �?              �?      .@              @              M@      (@       @      @               @       @       @       @      �?      �?      �?      �?                      �?      L@       @      B@       @      8@       @      &@       @      $@      �?      @      �?       @              @      �?      @              �?      �?      *@              (@              4@      @      (@      @      &@      �?      @      �?       @      �?              �?       @               @              @              �?      @              @      �?               @              A@      $@      @              =@      $@      @      "@               @      @      @      @       @       @      �?              �?       @              @      �?      �?      �?              �?      �?               @               @      @       @                      @      6@      �?      $@      �?      @      �?              �?      @              @              (@              D@      �?      0@      �?      @      �?      @                      �?      &@              8@              9@     �K@      @     �@@      @      (@      @      �?              �?      @                      &@              5@      4@      6@       @      1@              .@       @       @       @      �?      @              @      �?       @      �?      �?              �?      �?              �?      �?              �?                      �?      (@      @      $@               @      @              @       @      �?       @                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ��.hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM=huh*h-K ��h/��R�(KM=��h|�B@O         h                    �?��!h
��?�           @�@                                   �?N��6z�?�            �m@                                   �?���5��?$            �L@                                 �-@�T|n�q�?            �E@                                H�%@      �?             @        ������������������������       �                     �?        ������������������������       �                     @                                  �H@��-�=��?            �C@       	       
                   �;@г�wY;�?             A@        ������������������������       �        
             2@                                hf5@      �?             0@                                   �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        
             *@                                   �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        	             ,@               g                    @$�ݏ^��?p            �f@              *                     @�3_�4��?k            �e@                                  �?@�)�n�?7            @U@        ������������������������       �                     @                                    �?x�G�z�?4             T@                                  �:@�X�<ݺ?             B@                                   �?����X�?             @       ������������������������       �                     @                                  �8@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     =@                !                   @4@`���i��?             F@        ������������������������       �                     8@        "       #                    �?P���Q�?             4@        ������������������������       �                     @        $       )                    �?��S�ۿ?
             .@        %       &                    7@�q�q�?             @        ������������������������       �                     �?        '       (                    <@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     (@        +       f                 �̼6@�eP*L��?4             V@       ,       e                    @J�����?+            @S@       -       <                   �5@:W��S��?*             S@        .       /                    @����X�?             5@        ������������������������       �                      @        0       1                  s�@���y4F�?	             3@        ������������������������       �                     @        2       5                    �?����X�?             ,@        3       4                   �2@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        6       7                 @3"@"pc�
�?             &@        ������������������������       �                     @        8       9                    �?���Q��?             @        ������������������������       �                      @        :       ;                 ��l.@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        =       d                     @���Q��?            �K@       >       C                   �8@l`N���?            �J@        ?       B                   �7@؇���X�?             @       @       A                 ��Y@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        D       [                    �?(옄��?             G@       E       X                    �?     ��?             @@       F       M                    �?����"�?             =@        G       H                  ��@������?             .@        ������������������������       �                     �?        I       L                 �&B@d}h���?             ,@       J       K                 ���@�z�G��?             $@        ������������������������       �                     @        ������������������������       �և���X�?             @        ������������������������       �                     @        N       S                 ��� @      �?             ,@       O       R                   �;@�q�q�?             "@       P       Q                 �&B@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        T       U                    A@z�G�z�?             @        ������������������������       �                      @        V       W                    I@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        Y       Z                 ��"@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        \       ]                    .@և���X�?	             ,@        ������������������������       �                     @        ^       c                    �?      �?              @       _       `                    �?����X�?             @        ������������������������       �                     @        a       b                 ��1@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        	             &@        ������������������������       �                     @        i       �                    �?�՘���?'           �}@        j       k                 ���@R�����?1             T@        ������������������������       �                     @        l       �                    �?�;�vv��?+            @R@       m       �                  I>@��
ц��?              J@       n       �                   �=@b�2�tk�?             B@       o       |                 @Q,@l��[B��?             =@       p       q                     @�ՙ/�?	             5@        ������������������������       �                     �?        r       y                   @@���Q��?             4@       s       t                    5@��S���?             .@        ������������������������       �                     @        u       v                    9@�q�q�?             (@        ������������������������       �                     �?        w       x                   @<@�eP*L��?             &@       ������������������������       �      �?             $@        ������������������������       �                     �?        z       {                   �<@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        }       ~                   �8@      �?              @        ������������������������       �                     @               �                 `v�0@z�G�z�?             @        ������������������������       �                      @        �       �                    ;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                  �}S@      �?             0@       �       �                 �D�G@z�G�z�?             $@        �       �                 `f�A@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                 ��hU@�q�q�?             @        ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        �       �                   �H@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 �̾w@�ՙ/�?             5@       �       �                     �?��.k���?
             1@        �       �                   @K@      �?              @       ������������������������       �                     @        ������������������������       �                      @        �       �                   �6@�<ݚ�?             "@       �       �                    �?      �?              @        ������������������������       �                     @        �       �                 ��&@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �                          �?֓��H�?�            �x@       �       �                   �8@����?�             t@        �       �                   �3@��
���?/            �R@        �       �                    &@HP�s��?             9@       �       �                   �2@      �?             0@        ������������������������       �                      @        �       �                    �?      �?              @        ������������������������       �                     �?        �       �                 �?�@����X�?             @        ������������������������       �                     @        �       �                     @      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     I@        �       �                    �?V}�c
�?�            �n@        �       �                    �?�r����?             >@       �       �                   �=@ �Cc}�?             <@       �       �                   �:@؇���X�?             5@        ������������������������       �                     �?        �       �                    �?R���Q�?             4@       �       �                 `ff@z�G�z�?	             .@        ������������������������       �                     @        ������������������������       ����!pc�?             &@        ������������������������       �                     @        ������������������������       �                     @        �       �                    B@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �;@�*�����?�             k@        �       �                   �:@     ��?             @@       �       �                     @���N8�?             5@        ������������������������       �                     @        �       �                 `�B@�q�q�?             .@       �       �                   �9@�θ�?
             *@        �       �                 @33@և���X�?             @        ������������������������       �                     �?        �       �                    �?�q�q�?             @        ������������������������       �                     @        �       �                 (3�)@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                     �?�C��2(�?             &@        ������������������������       �                     @        �       �                 ��T1@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                     �?t��eh��?y             g@        �       �                   @I@�+e�X�?             I@       �       �                    D@r�q��?             E@       �       �                   �B@�θ�?             :@       �       �                   �A@z�G�z�?             9@       �       �                 ��yC@��<b���?             7@       �       �                 ��$:@X�Cc�?
             ,@        ������������������������       �                     @        �       �                   �?@      �?              @       �       �                 `fF<@և���X�?             @        ������������������������       �                     �?        �       �                   �>@�q�q�?             @        ������������������������       �                     @        �       �                   �A@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?      �?             0@       �       �                 `f�;@�C��2(�?             &@       �       �                 ��:@      �?             @        ������������������������       �                     �?        �       �                   @G@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   �J@      �?              @        ������������������������       �                     @        �       �                   �Q@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                 �?�@\��ut-�?[            �`@        �       �                 ���@�(\����?             D@        ������������������������       �                     2@        �       �                 �?$@���7�?             6@        �       �                   �>@      �?             @        ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     2@        �                          �?�!��U��?>            �W@       �                        @3�@���y4F�?0             S@        �       �                    C@����X�?             @       �       �                   �?@���Q��?             @        ������������������������       �                     �?        ������������������������       �      �?             @        ������������������������       �                      @                                @@@0)RH'�?,            @Q@                             ��y @�θ�?            �C@                              ��) @ҳ�wY;�?
             1@                                ?@8�Z$���?	             *@       ������������������������       �                     &@        ������������������������       �                      @        ������������������������       �                     @                                @<@��2(&�?             6@       	                          @z�G�z�?             .@        
                        �*@���Q��?             @                               �'@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @                              �T�C@ףp=
�?             $@       ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                     @                                `M@��S�ۿ?             >@                               @A@h�����?             <@                                �@@�����H�?             "@        ������������������������       �                     @                              ��%@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     3@                                �P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     3@                                  �?X~�pX��?)            @R@        ������������������������       �                     @        !      0                    @.Lj���?&             Q@        "      +                 x�N@`՟�G��?             ?@       #      $                   �?������?
             1@        ������������������������       �                      @        %      &                    �?�r����?	             .@        ������������������������       �                     @        '      (                   :@"pc�
�?             &@        ������������������������       �                     @        )      *                  �9@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ,      /                   �?@4և���?             ,@        -      .                   )@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        1      <                   @���"͏�?            �B@       2      ;                   @�z�G��?             >@       3      6                   �?     ��?	             0@       4      5                    @�eP*L��?             &@        ������������������������       �                     @        ������������������������       �                     @        7      8                ���9@z�G�z�?             @        ������������������������       �                      @        9      :                ��T?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     ,@        ������������������������       �                     @        �t�bh�h*h-K ��h/��R�(KM=KK��h]�B�       �z@     �q@     @P@     �e@      @      I@      @      B@      @      �?              �?      @              @     �A@      �?     �@@              2@      �?      .@      �?       @               @      �?                      *@      @       @      @                       @              ,@      M@     �^@     �I@     �^@      @     �T@              @      @     @S@       @      A@       @      @              @       @      �?              �?       @                      =@      �?     �E@              8@      �?      3@              @      �?      ,@      �?       @              �?      �?      �?      �?                      �?              (@      H@      D@     �B@      D@     �B@     �C@      .@      @               @      .@      @      @              $@      @      �?       @               @      �?              "@       @      @              @       @       @              �?       @               @      �?              6@     �@@      6@      ?@      �?      @      �?       @               @      �?                      @      5@      9@      *@      3@      &@      2@      @      &@      �?              @      &@      @      @              @      @      @              @      @      @      @      @      �?      @      �?                      @      @              �?      @               @      �?       @      �?                       @       @      �?       @                      �?       @      @      @               @      @       @      @              @       @      �?              �?       @                      �?               @              �?      &@              @             �v@     �[@     �E@     �B@      @              B@     �B@      <@      8@      6@      ,@      .@      ,@       @      *@              �?       @      (@      @       @              @      @      @      �?              @      @      @      @      �?              �?      @      �?                      @      @      �?      @              @      �?       @               @      �?              �?       @              @              @      $@       @       @       @      @              @       @                      @      @       @      @              �?       @              �?      �?      �?              �?      �?               @      *@       @      "@      @       @      @                       @       @      @      �?      @              @      �?      @      �?                      @      �?                      @      t@     @R@      q@      I@     @R@       @      7@       @      ,@       @       @              @       @      �?              @       @      @               @       @       @      �?              �?      "@              I@             �h@      H@      :@      @      9@      @      2@      @      �?              1@      @      (@      @      @               @      @      @              @              �?      �?              �?      �?             �e@      F@      1@      .@      0@      @      @              $@      @      $@      @      @      @              �?      @       @      @              �?       @               @      �?              @                       @      �?      $@              @      �?      @              @      �?             �c@      =@      C@      (@     �A@      @      4@      @      4@      @      2@      @      "@      @      @              @      @      @      @      �?               @      @              @       @      �?       @                      �?              �?      "@               @                      �?      .@      �?      $@      �?      @      �?      �?               @      �?       @                      �?      @              @              @      @              @      @       @      @                       @     �]@      1@     �C@      �?      2@              5@      �?      @      �?      �?      �?       @              2@             �S@      0@      N@      0@       @      @       @      @              �?       @       @               @      M@      &@      >@      "@      &@      @      &@       @      &@                       @              @      3@      @      (@      @      @       @      �?       @      �?                       @       @              "@      �?      @               @      �?      @              <@       @      ;@      �?       @      �?      @               @      �?       @                      �?      3@              �?      �?              �?      �?              3@              I@      7@      @             �F@      7@      1@      ,@      @      *@       @               @      *@              @       @      "@              @       @      @              @       @              *@      �?      @      �?              �?      @              @              <@      "@      5@      "@      @      "@      @      @              @      @              �?      @               @      �?       @      �?                       @      ,@              @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJj�c;hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM-huh*h-K ��h/��R�(KM-��h|�B@K         ^                    �?�)�>_M�?�           @�@               M                    �?�T����?�            0p@                                  �?�����?�            �l@                                   �?�t����?5            @U@              
                     @�F��O�?.            @R@                                 �H@�Ń��̧?             E@       ������������������������       �                     A@               	                 83F@      �?              @        ������������������������       �                     �?        ������������������������       �                     @                                   �?�חF�P�?             ?@                                   7@���!pc�?             &@                               P��+@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @                                   7@ףp=
�?             4@                                 s�@      �?             @        ������������������������       �                     �?        ������������������������       �                     @                                   �?      �?	             0@                               pF @ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     @                                ���.@�q�q�?             (@        ������������������������       �                     @        ������������������������       �                      @               *                     @�ň?�S�?Z             b@                                  @��+��<�?6            �U@        ������������������������       �                     �?                )                   �;@�D�e���?5            @U@        !       "                   �8@ 	��p�?             =@       ������������������������       �                     7@        #       &                    :@�q�q�?             @       $       %                     �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        '       (                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        #             L@        +       ,                 ���@�Ƀ aA�?$            �M@        ������������������������       �                      @        -       F                    �?�q�q�?             �I@       .       ;                    �?�ՙ/�?             E@       /       4                 ��&@������?             >@       0       3                    3@P���Q�?             4@        1       2                 x&�!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        
             2@        5       :                 03�1@�z�G��?             $@       6       9                 ��Y.@      �?              @        7       8                 ���*@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        <       E                 0336@�q�q�?             (@       =       B                    <@z�G�z�?             $@       >       A                 P��%@      �?              @        ?       @                   �#@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        C       D                    @@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        G       L                    �?�����H�?             "@        H       K                    @      �?             @       I       J                    @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        N       U                    �?����"�?             =@        O       T                    @����X�?             @       P       Q                      @      �?             @        ������������������������       �                     �?        R       S                    7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        V       ]                 ���d@���!pc�?             6@       W       X                    @�IєX�?             1@        ������������������������       �                     $@        Y       \                    @؇���X�?             @        Z       [                 ��T?@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        _       t                    $@�g[Z��?            P|@        `       i                    �?և���X�?             <@       a       h                    !@X�<ݚ�?             2@       b       c                   �;@և���X�?
             ,@        ������������������������       �                     @        d       e                   A@�����H�?             "@       ������������������������       �                     @        f       g                   �C@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        j       k                    �?���Q��?             $@        ������������������������       �                      @        l       s                  DP@      �?              @       m       r                    @�q�q�?             @       n       o                 ���9@�q�q�?             @        ������������������������       �                     �?        p       q                 ��T?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        u       �                    �?���f_�?           �z@        v       �                 83##@�	j*D�?2            �S@        w       z                    5@�C��2(�?            �@@        x       y                 �{@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        {       �                    =@`Jj��?             ?@       |       }                 ���@ףp=
�?             4@        ������������������������       �                     @        ~                           9@؇���X�?             ,@        ������������������������       �                      @        �       �                   @@r�q��?             (@       ������������������������       �z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                     &@        �       �                    �?��S���?            �F@       �       �                    I@X��ʑ��?            �E@       �       �                    �?��
ц��?            �C@       �       �                   �8@�eP*L��?             6@        �       �                     �?      �?             @        �       �                   �3@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �;@b�2�tk�?             2@        ������������������������       �                     @        �       �                 �;|r@��S���?
             .@       �       �                    A@��
ц��?	             *@       �       �                     �?���Q��?             $@       �       �                    ?@X�<ݚ�?             "@       �       �                 ���<@և���X�?             @       ������������������������       �                     @        �       �                 03SA@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    D@��.k���?             1@       �       �                     @�n_Y�K�?	             *@       �       �                   �:@�<ݚ�?             "@        �       �                     �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?      �?             @       �       �                    3@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �                       ��$:@�-q���?�            �u@       �       �                    �?dP-���?�            �q@       �       �                     �?��(\���?�             n@        ������������������������       �                     $@        �       �                    1@ج��w�?�            �l@        �       �                     @      �?              @        ������������������������       �                      @        �       �                 pFD!@      �?             @        �       �                 pf�@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                 ���"@,N�_� �?�            �k@       �       �                   �@���	���?_            �b@       �       �                  ��@�L���?2            �R@       �       �                   �;@ �#�Ѵ�?            �E@        �       �                    �?      �?             0@        ������������������������       �                      @        �       �                 ���@؇���X�?	             ,@       �       �                    :@�<ݚ�?             "@       �       �                 ���@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     ;@        �       �                    �?��� ��?             ?@        �       �                   �>@r�q��?	             (@       �       �                 ��(@�<ݚ�?             "@       �       �                   �<@����X�?             @       ������������������������       �r�q��?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                 �?$@�KM�]�?             3@        ������������������������       �                      @        �       �                 �1@"pc�
�?             &@        �       �                   �6@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 P�N@؇���X�?             @        ������������������������       �                     �?        �       �                   �:@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    ?@�e���@�?-            @S@       ������������������������       �        "            �N@        �       �                 @3�@      �?             0@        ������������������������       �                     @        �       �                   �@@ףp=
�?             $@        �       �                 ��i @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                     @�Z��L��?*            �Q@       �       �                   @N@��2(&�?             F@       �       �                   �*@X�EQ]N�?            �E@       �       �                 `f�)@�>4և��?             <@        ������������������������       �                     "@        �       �                    C@�d�����?             3@       �       �                    =@ףp=
�?             $@        �       �                    :@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �F@X�<ݚ�?             "@        ������������������������       �z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     .@        ������������������������       �                     �?        �       �                   �<@�>����?             ;@       ������������������������       �                     .@        �       �                    �?r�q��?             (@       �       �                 03�0@����X�?             @       �       �                    ?@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �                         �9@؇���X�?             E@        �                       pf(@X�Cc�?	             ,@       �                          �?X�<ݚ�?             "@       �                          �7@      �?              @       �       �                 ��Y@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @                                 �?h�����?             <@       ������������������������       �                     4@                                 �?      �?              @                                ;@؇���X�?             @        ������������������������       �                     @        	      
                   �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?              $                    �?؇>���?-            @P@                               �>@������?            �D@                                 L@և���X�?             ,@                               `G@z�G�z�?
             $@                               �F@      �?              @                               �?@؇���X�?             @                             `fF<@      �?             @        ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @              #                  �C@PN��T'�?             ;@                               �=@������?
             1@       ������������������������       �                      @                                 �@@X�<ݚ�?             "@                                @K@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        !      "                03�X@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        	             $@        %      ,                   �?r�q��?             8@        &      +                ��?P@����X�?             ,@       '      *                   >@      �?              @       (      )                   ;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �z�G�z�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     $@        �t�bh�h*h-K ��h/��R�(KM-KK��h]�B�       `{@      q@     @P@     @h@     �G@     �f@      $@     �R@      @     �P@      �?     �D@              A@      �?      @      �?                      @      @      :@      @       @      @      @              @      @                      @       @      2@      �?      @      �?                      @      �?      .@      �?      "@              "@      �?                      @      @       @      @                       @     �B@      [@      @     �T@      �?               @     �T@       @      ;@              7@       @      @      �?       @      �?                       @      �?       @               @      �?                      L@      A@      9@               @      A@      1@      :@      0@      6@       @      3@      �?      �?      �?      �?                      �?      2@              @      @      �?      @      �?       @               @      �?                      @       @              @       @       @       @      �?      @      �?      �?              �?      �?                      @      �?      �?      �?                      �?       @               @      �?      @      �?       @      �?              �?       @              �?              @              2@      &@       @      @       @       @              �?       @      �?       @                      �?              @      0@      @      0@      �?      $@              @      �?       @      �?       @                      �?      @                      @     Pw@      T@      (@      0@       @      $@       @      @              @       @      �?      @               @      �?              �?       @                      @      @      @               @      @      @      @       @      �?       @              �?      �?      �?      �?                      �?      @                       @     �v@      P@      K@      8@      >@      @      �?      �?      �?                      �?      =@       @      2@       @      @              (@       @       @              $@       @       @       @       @              &@              8@      5@      6@      5@      2@      5@      $@      (@      @      �?      �?      �?              �?      �?               @              @      &@              @      @       @      @      @      @      @      @      @      @      @      @              �?      @              @      �?                       @              �?      @                       @       @      "@       @      @      @       @       @       @               @       @              @              �?      @      �?      �?              �?      �?                       @              @      @               @             0s@      D@      p@      8@     �k@      2@      $@             �j@      2@      @      @       @              @      @      �?      @      �?                      @       @             �i@      .@      b@      @      Q@      @     �D@       @      ,@       @       @              (@       @      @       @      @      �?      @                      �?              �?      @              ;@              ;@      @      $@       @      @       @      @       @      @      �?              �?       @              @              1@       @       @              "@       @      @      �?              �?      @              @      �?      �?              @      �?      @                      �?      S@      �?     �N@              .@      �?      @              "@      �?       @      �?              �?       @              @             �O@       @      C@      @      C@      @      7@      @      "@              ,@      @      "@      �?      @      �?      @                      �?      @              @      @      �?      @      @              .@                      �?      9@       @      .@              $@       @      @       @      @       @               @      @               @              @              B@      @      "@      @      @      @      @      @      @       @      @                       @              @      �?              @              ;@      �?      4@              @      �?      @      �?      @              @      �?              �?      @              �?             �H@      0@      =@      (@      @       @       @       @       @      @      �?      @      �?      @      �?      �?               @              @      �?                       @      @              7@      @      *@      @       @              @      @      @       @      @                       @       @       @       @                       @      $@              4@      @      $@      @      @      @      @       @              �?      @      �?               @      @              $@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJGԙGhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM[huh*h-K ��h/��R�(KM[��h|�B�V         �                     @�3�n��?�           @�@                                  �'@z�J��?�            �t@                                   �?      �?             D@        ������������������������       �                     @                                    �?@-�_ .�?            �B@        ������������������������       �                     @                                  �H@��S�ۿ?             >@              	                    @ 7���B�?             ;@        ������������������������       �                      @        
                           4@�}�+r��?
             3@                                  �2@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     (@                                  �P@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @               {                   �J@D$f�y�?�            r@              z                    �?      �?x             h@                                 �6@�Ҵ$��?t            `g@                                   �?���}<S�?             7@       ������������������������       �        	             1@                                   �?�q�q�?             @        ������������������������       �                     �?                                  `?@z�G�z�?             @        ������������������������       �                     @                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               9                 �̌-@yÏP�?f            �d@               "                    �?H(���o�?            �J@                !                   �E@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        #       8                    �?���Q��?            �F@       $       )                    �?8�A�0��?             F@        %       &                 `f�)@���}<S�?
             7@        ������������������������       �                     @        '       (                    :@�����H�?	             2@        ������������������������       ��q�q�?             @        ������������������������       �                     (@        *       7                   �*@���N8�?             5@       +       ,                   �:@�t����?             1@        ������������������������       �                     @        -       .                    =@�q�q�?             (@        ������������������������       �                     @        /       0                 `f�)@�<ݚ�?             "@        ������������������������       �                     �?        1       2                    @@      �?              @        ������������������������       �                     �?        3       4                   @B@����X�?             @        ������������������������       �      �?              @        5       6                   @D@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     �?        :       E                    �?4�B��?H            �[@        ;       >                    �?�C��2(�?             6@        <       =                   �H@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ?       @                    �?�}�+r��?             3@        ������������������������       �                      @        A       D                    <@�C��2(�?             &@        B       C                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        F       s                   @H@&<k����?8            @V@       G       r                    �?� ���?.            @S@       H       S                 ��$:@"pc�
�?'            �P@        I       J                    9@ 7���B�?             ;@        ������������������������       �                     &@        K       L                     �?      �?	             0@        ������������������������       �                      @        M       N                    �?@4և���?             ,@        ������������������������       �                     @        O       R                   �@@؇���X�?             @        P       Q                   �<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        T       U                   �;@�(�Tw��?            �C@        ������������������������       �                     �?        V       _                    �?�d�����?             C@        W       ^                 `f�A@      �?              @       X       ]                   �>@���Q��?             @       Y       \                     �?�q�q�?             @       Z       [                 �ܵ<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        `       q                     �?�������?             >@       a       b                 03k:@>���Rp�?             =@        ������������������������       �                     @        c       p                 ��yC@8�Z$���?             :@       d       i                   @=@�	j*D�?	             *@        e       h                 `f�;@z�G�z�?             @       f       g                   @B@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     �?        j       o                   �<@      �?              @       k       l                   @@@      �?             @        ������������������������       �                      @        m       n                   �A@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     *@        ������������������������       �                     �?        ������������������������       �                     &@        t       u                    �?�q�q�?
             (@        ������������������������       �                     �?        v       y                    @@���!pc�?	             &@       w       x                   �J@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        |       �                    �?�^�X�?C            @X@       }       �                    �?@�h�|5�?=            @V@       ~                         "�b@h㱪��?$            �K@       ������������������������       �                    �D@        �       �                    �?؇���X�?
             ,@       ������������������������       �                     &@        �       �                    <@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?ҳ�wY;�?             A@       �       �                    �?��S���?             .@       �       �                   �7@�eP*L��?	             &@        ������������������������       �                     @        �       �                  �}S@      �?              @        ������������������������       �                     @        �       �                 0�HU@      �?             @        ������������������������       �                     �?        �       �                    �?�q�q�?             @       �       �                   �?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   PP@      �?             @        ������������������������       �                     �?        �       �                   �B@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?���y4F�?             3@       �       �                    �?�q�q�?             "@        �       �                   �4@�q�q�?             @        ������������������������       �                     �?        �       �                    >@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 `��S@r�q��?             @        ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                ����8@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        �       �                    �?      �?              @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�E�_�?�            �w@        �       �                    �?؇���X�?             @       ������������������������       �                     @        �       �                 8#8@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?@�҇��?�            �w@        �       �                   �>@$ޗQ��?A            �Y@       �       �                 03�7@ 9�����?8             V@       �       �                    �?a��t��?3            �S@       �       �                    �?D������?,            @P@        �       �                    �?����e��?            �@@        �       �                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?l��
I��?             ;@       �       �                    �?`�Q��?             9@       �       �                   �<@�q�q�?             8@       �       �                    ;@�GN�z�?             6@        �       �                   �9@���Q��?             @       �       �                   �0@�q�q�?             @        ������������������������       �                     �?        �       �                   �7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ���@�t����?
             1@        ������������������������       �                     @        �       �                   @<@"pc�
�?             &@       �       �                   @@z�G�z�?             $@       ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �5@     ��?             @@        �       �                    �?z�G�z�?             @       �       �                   �0@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?��}*_��?             ;@       �       �                    �?���Q��?             9@       �       �                  ��@���|���?             6@        ������������������������       �                      @        �       �                    9@�z�G��?             4@        ������������������������       �                     �?        �       �                    �?�����?             3@       �       �                 pF @     ��?
             0@       �       �                 �&B@@4և���?	             ,@       �       �                 ���@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �ףp=
�?             $@        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                 ���.@�θ�?             *@       �       �                    �?      �?             @        �       �                 P��+@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �<@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �        	             ,@        �       &                   �?����c�?�             q@        �                       ���4@���3E��?8            @W@       �                          @     8�?&             P@       �                         �9@V{q֛w�?%             O@        �                          �?��>4և�?             <@       �       �                 ���@��}*_��?             ;@        ������������������������       �                     @        �                          �?�GN�z�?             6@       �       �                  �#@@�0�!��?	             1@       ������������������������       �                     &@        �       �                    �?      �?             @        �       �                    4@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �                          �&@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                              �̬)@���Q��?             @        ������������������������       �                      @                                 �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?                                �;@�t����?             A@        	                        �:@$�q-�?             *@        
                         �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @                                 =@և���X�?             5@                                 �?����X�?             @                                �?�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?                                 �?����X�?	             ,@                               @B@�q�q�?             (@                             03�1@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?                                 �?���Q��?             @                                I@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @               !                   �?XB���?             =@        ������������������������       �                      @        "      %                   @���N8�?             5@        #      $                   @      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     1@        '      Z                   �?�����?s            �f@       (      Y                   �?���Ehz�?h            �d@       )      *                   $@\���(�?d             d@        ������������������������       �                     �?        +      R                   �?�NW���?c            �c@       ,      O                �T�C@ȥ�fzR�?S             a@       -      .                �&B@P�2E��?O            @`@        ������������������������       �                     B@        /      4                �{@=QcG��?:            �W@        0      1                  �:@����X�?             @        ������������������������       �                     @        2      3                   D@      �?             @        ������������������������       �                      @        ������������������������       �                      @        5      8                  �0@`��F:u�?7            �U@        6      7                pFD!@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        9      B                   ?@h�����?5             U@       :      ;                  �:@     ��?%             P@       ������������������������       �                     A@        <      =                pf� @(;L]n�?             >@       ������������������������       �                     4@        >      A                ��)"@ףp=
�?             $@        ?      @                  �;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        C      H                  @@@ףp=
�?             4@        D      E                @3�@z�G�z�?             @        ������������������������       �                     @        F      G                ��i @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        I      J                  �E@��S�ۿ?             .@        ������������������������       �                      @        K      N                  �F@؇���X�?             @        L      M                @3�@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        P      Q                   ;@և���X�?             @        ������������������������       �                      @        ������������������������       ����Q��?             @        S      X                  �9@�C��2(�?             6@        T      U                ��@r�q��?             (@        ������������������������       �                     @        V      W                �&B@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                     @        ������������������������       �                     .@        �t�b��2     h�h*h-K ��h/��R�(KM[KK��h]�B�       �{@     �p@      d@      e@     �A@      @              @     �A@       @      @              <@       @      :@      �?       @              2@      �?      @      �?      @                      �?      (@               @      �?              �?       @             �_@     `d@      X@      X@      X@     �V@       @      5@              1@       @      @      �?              �?      @              @      �?      �?              �?      �?             �W@     �Q@      3@      A@      �?      @              @      �?              2@      ;@      2@      :@       @      5@              @       @      0@       @      @              (@      0@      @      (@      @      @              @      @              @      @       @      �?              @       @      �?              @       @      �?      �?      @      �?      �?              @      �?      @                      �?     �R@      B@       @      4@      �?       @               @      �?              �?      2@               @      �?      $@      �?      @      �?                      @              @     @R@      0@     @P@      (@      K@      (@      :@      �?      &@              .@      �?       @              *@      �?      @              @      �?      �?      �?      �?                      �?      @              <@      &@              �?      <@      $@      @      @       @      @       @      �?      �?      �?      �?                      �?      �?                       @      @              7@      @      6@      @              @      6@      @      "@      @      @      �?      @      �?      �?               @      �?      �?              @      @      �?      @               @      �?      �?      �?                      �?      @              *@              �?              &@               @      @              �?       @      @      @      @              @      @              @                      @      >@     �P@      8@     @P@       @     �J@             �D@       @      (@              &@       @      �?       @                      �?      6@      (@      @       @      @      @      @               @      @              @       @       @      �?              �?       @      �?      �?      �?                      �?              �?       @       @              �?       @      �?       @                      �?      .@      @      @      @      �?       @              �?      �?      �?      �?                      �?      @      �?      @              �?      �?      �?                      �?      "@      �?              �?      "@              @       @               @      @             �q@     �X@      �?      @              @      �?      �?              �?      �?             �q@      W@     �N@     �D@     �G@     �D@     �B@     �D@      A@      ?@      4@      *@      �?      @              @      �?              3@       @      1@       @      1@      @      1@      @       @      @       @      �?      �?              �?      �?              �?      �?                       @      .@       @      @              "@       @       @       @      @       @       @              �?                       @              �?       @              ,@      2@      @      �?       @      �?              �?       @               @              $@      1@      $@      .@       @      ,@       @              @      ,@              �?      @      *@      @      *@      �?      *@      �?      $@              �?      �?      "@              @       @              @               @      �?              �?       @                       @      @      $@      @      @      �?      �?              �?      �?               @       @       @                       @              @      $@              ,@             �k@     �I@     �K@      C@      ;@     �B@      ;@     �A@      1@      &@      1@      $@              @      1@      @      ,@      @      &@              @      @       @       @               @       @              �?      �?      �?                      �?      @       @       @              �?       @               @      �?                      �?      $@      8@      �?      (@      �?      @              @      �?                      @      "@      (@      @       @      @       @      @                       @      �?              @      $@      @       @      �?      @              @      �?              @       @       @       @       @                       @      �?                       @               @      <@      �?       @              4@      �?      @      �?      @                      �?      1@              e@      *@      c@      *@     `b@      *@              �?     `b@      (@     �_@      $@      _@      @      B@              V@      @      @       @      @               @       @               @       @             �T@      @       @      �?              �?       @             @T@      @     �O@      �?      A@              =@      �?      4@              "@      �?      �?      �?              �?      �?               @              2@       @      @      �?      @              �?      �?              �?      �?              ,@      �?       @              @      �?      �?      �?              �?      �?              @              @      @               @      @       @      4@       @      $@       @      @              @       @               @      @              $@              @              .@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ��AhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM7huh*h-K ��h/��R�(KM7��h|�B�M         b                    �?ƈ�VM�?�           @�@               a                    @2�K^V�?�            �p@              Z                   XB@ja_e���?�            pp@                                   @Fe5]�>�?p            `f@               
                     �?h�����?'             L@                                `v7<@����X�?             @       ������������������������       �                     @               	                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        "            �H@               U                 `v�6@.M�d�c�?I            �^@              (                    �?�$q�Y	�??            @[@                                  �+@>��C��?            �E@        ������������������������       �                     $@               #                    �?:ɨ��?            �@@              "                    �?`�Q��?             9@                                  �?�GN�z�?             6@                                   0@z�G�z�?             @        ������������������������       �                      @                                  �6@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                  �8@������?             1@                                  �0@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                ���@؇���X�?             ,@        ������������������������       �                     �?                                 s�@$�q-�?             *@        ������������������������       �                     @                !                 �&B@ףp=
�?             $@       ������������������������       �؇���X�?             @        ������������������������       �                     @        ������������������������       �                     @        $       '                    �?      �?              @       %       &                    �?����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        )       H                    �?�\����?'            �P@       *       G                    A@�~8�e�?            �I@       +       F                    �?      �?             F@       ,       ?                   �:@�G��l��?             E@       -       :                    �?*;L]n�?             >@       .       /                 ���@�eP*L��?             6@        ������������������������       �                     "@        0       9                 pf� @�θ�?
             *@       1       6                 P�@      �?              @       2       3                    4@z�G�z�?             @        ������������������������       �                     @        4       5                   �7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        7       8                   �8@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ;       <                 �̬)@      �?              @       ������������������������       �                     @        =       >                 @3�/@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        @       E                    �?      �?             (@       A       D                 ��� @և���X�?             @       B       C                   �;@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        I       T                    @�r����?
             .@       J       S                    �?8�Z$���?	             *@       K       N                    $@z�G�z�?             $@        L       M                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        O       P                   �*@      �?              @        ������������������������       �                     @        Q       R                 03S1@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        V       W                 ��T?@؇���X�?
             ,@       ������������������������       �                     "@        X       Y                    @���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        [       \                 ���a@�Ń��̧?5             U@       ������������������������       �        (             N@        ]       ^                    !@�8��8��?             8@        ������������������������       �                     �?        _       `                 03c@�nkK�?             7@        ������������������������       �                     �?        ������������������������       �                     6@        ������������������������       �                      @        c                       `fFJ@�����?           �{@       d       {                    �?�=�w\�?�             x@        e       z                    �?�I�w�"�?             C@       f       u                 ���<@<���D�?            �@@       g       t                    �?ܷ��?��?             =@       h       k                     @�����H�?             ;@        i       j                     �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        l       o                   �7@���}<S�?             7@        m       n                    5@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        p       s                   @<@�X�<ݺ?             2@       q       r                 ���@�C��2(�?             &@        ������������������������       �                     @        ������������������������       �r�q��?             @        ������������������������       �                     @        ������������������������       �                      @        v       y                    @@      �?             @       w       x                 03SA@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        |       �                     �?r�q��?�            �u@        }       �                    �?�+e�X�?             I@       ~       �                   �>@��+7��?             G@              �                 `fF<@
j*D>�?             :@       �       �                 ��$:@������?
             1@        ������������������������       �                     @        �       �                 03k:@���Q��?             $@        ������������������������       �                     �?        �       �                    K@�q�q�?             "@        �       �                    C@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   �<@�<ݚ�?             "@        ������������������������       �                     @        �       �                   �P@      �?             @       ������������������������       �                      @        ������������������������       �                      @        �       �                   �=@P���Q�?
             4@        �       �                   �A@ףp=
�?             $@        ������������������������       �                     @        �       �                 ��yC@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �                     @        �       �                 �?�@,:#\��?�            �r@        �       �                    �?d����?D            �\@        �       �                  ��@      �?             4@        ������������������������       �                     @        �       �                   �<@X�Cc�?             ,@       �       �                 ��(@�<ݚ�?             "@       ������������������������       �      �?              @        ������������������������       �                     �?        �       �                   �>@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                     @<����?9            �W@        ������������������������       �                     @        �       �                    �?�:�^���?6            �V@       �       �                 ��@�^;\��?5            @V@        �       �                 @3�@      �?             $@        �       �                   �B@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �>@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �@(�5�f��?/            �S@       �       �                 �?$@��<D�m�?            �H@       �       �                   �8@P�Lt�<�?             C@        �       �                    7@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     >@        �       �                 ��L@"pc�
�?             &@        �       �                   �5@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �:@؇���X�?             @        ������������������������       �                     @        �       �                    D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     >@        ������������������������       �                     �?        �       �                 @3�@L=�m��?v            �f@        �       �                    :@և���X�?             @        ������������������������       �                     �?        �       �                    �?      �?             @       �       �                   �?@���Q��?             @        ������������������������       �                     �?        ������������������������       �      �?             @        ������������������������       �                     �?        �       �                    @��!pc�?p             f@        �       �                     @d}h���?	             ,@       ������������������������       �                      @        �       �                 ��|2@      �?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                 ��y)@����ր�?g            @d@        �       �                    &@z��R[�?/            �Q@        ������������������������       �                      @        �       �                    �?�� =[�?-             Q@       �       �                   �=@� y���?,            �P@       �       �                 ���!@H.�!���?"             I@       �       �                 ��) @�q�q�?             8@       �       �                    4@      �?             0@        �       �                   �1@z�G�z�?             @       ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �        
             &@        �       �                 pf� @      �?              @        ������������������������       �                     �?        �       �                    8@և���X�?             @       ������������������������       �                     @        �       �                   �;@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                 ���#@ȵHPS!�?             :@       �       �                   �<@@�0�!��?	             1@       ������������������������       �                     *@        �       �                 ���"@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �        
             1@        ������������������������       �                     �?        �       �                    �?���.�6�?8             W@        �       �                    2@�8��8��?             (@        ������������������������       �                     @        �       �                    A@r�q��?             @       �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �                          �?      �?1             T@       �                           �?�ӖF2��?+            �Q@       �       �                   @A@`Ӹ����?            �F@       �       �                     @�>����?             ;@       �       �                    �?�����H�?
             2@       �       �                   �3@      �?	             0@       �       �                   �:@�r����?             .@        ������������������������       �                     @        �       �                    =@�<ݚ�?             "@        ������������������������       �                     �?        �       �                    @@      �?              @        ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     2@                                 �?ȵHPS!�?             :@                                �?@�0�!��?             1@              
                    @      �?              @                               �<@r�q��?             @        ������������������������       �                     @              	                  �:@�q�q�?             @                               �@@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @                                  @�<ݚ�?             "@                                +@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @                              `f4@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     "@                              ��#@<|ۤ$�?!            �K@        ������������������������       �                      @              4                   �?Fmq��?             �J@             /                   �?X�<ݚ�?            �F@             .                     @�eP*L��?            �@@             %                   �?���>4��?             <@                                �?@j���� �?             1@                                �?���Q��?             $@        ������������������������       �                     @                                �:@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        !      "                @�pX@؇���X�?             @        ������������������������       �                     @        #      $                  @E@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        &      -                03�M@���!pc�?             &@       '      ,                ��9L@և���X�?             @       (      +                  @K@�q�q�?             @       )      *                   7@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        0      3                   �?r�q��?             (@       1      2                   L@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                     �?        5      6                  �G@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        �t�bh�h*h-K ��h/��R�(KM7KK��h]�Bp        z@     �r@     @P@     �i@     �L@     �i@     �K@      _@       @      K@       @      @              @       @      �?       @                      �?             �H@     �J@     �Q@     �D@      Q@      $@     �@@              $@      $@      7@       @      1@      @      1@      �?      @               @      �?       @      �?                       @      @      *@       @      �?              �?       @               @      (@      �?              �?      (@              @      �?      "@      �?      @              @      @               @      @       @      @       @                      @              �?      ?@     �A@      =@      6@      6@      6@      4@      6@      1@      *@      $@      (@              "@      $@      @      @      @      @      �?      @              �?      �?              �?      �?              �?       @      �?                       @      @              @      �?      @              @      �?              �?      @              @      "@      @      @      @       @               @      @                       @              @       @              @               @      *@       @      &@       @       @      �?      �?      �?                      �?      �?      @              @      �?      @      �?                      @              @               @      (@       @      "@              @       @               @      @               @     �T@              N@       @      6@      �?              �?      6@      �?                      6@       @             �u@     �V@     �s@     �P@      =@      "@      =@      @      :@      @      8@      @      @      �?      @                      �?      5@       @      @      �?      @                      �?      1@      �?      $@      �?      @              @      �?      @               @              @      �?      �?      �?              �?      �?               @                      @      r@      M@      C@      (@      A@      (@      .@      &@      *@      @      @              @      @              �?      @      @      �?      @      �?                      @      @               @      @              @       @       @       @                       @      3@      �?      "@      �?      @               @      �?              �?       @              $@              @             �o@      G@     �Y@      *@      .@      @      @              "@      @      @       @      @       @      �?               @      @              @       @             �U@       @      @             �T@       @     @T@       @      @      @      �?       @               @      �?              @      @              @      @              S@      @      G@      @     �B@      �?      @      �?      @                      �?      >@              "@       @      @      �?              �?      @              @      �?      @              �?      �?              �?      �?              >@              �?             �b@     �@@      @      @      �?              @      @       @      @              �?       @       @      �?             @b@      >@      @      &@               @      @      @              @      @             �a@      3@     �L@      *@               @     �L@      &@      L@      &@     �C@      &@      0@       @      (@      @      �?      @      �?       @               @      &@              @      @              �?      @      @      @              �?      @              @      �?              7@      @      ,@      @      *@              �?      @      �?                      @      "@              1@              �?             �U@      @      &@      �?      @              @      �?      @      �?      @                      �?       @             �R@      @     �P@      @     �E@       @      9@       @      0@       @      ,@       @      *@       @      @              @       @              �?      @      �?      @               @      �?      �?               @              "@              2@              7@      @      ,@      @      @      �?      @      �?      @               @      �?      �?      �?              �?      �?              �?               @              @       @      @      �?              �?      @              �?      �?              �?      �?              "@              "@              @@      7@               @      @@      5@      9@      4@      .@      2@      .@      *@      @      $@      @      @      @               @      @              @       @              �?      @              @      �?      @              @      �?               @      @      @      @      @       @       @       @       @                       @       @                      �?      @                      @      $@       @      $@      �?      $@                      �?              �?      @      �?      @                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ,�hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMQhuh*h-K ��h/��R�(KMQ��h|�B@T         �                     @\H�l�?�           @�@               Q                     �?d�2�,��?�            �r@               P                    @��g�ao�?[            �a@                                  �?nIz~]�?Z            �a@                                   "@$�q-�?&            @P@        ������������������������       �                     �?                                 "�b@      �?%             P@                                  �?�O4R���?            �J@       	                        03[=@      �?             @@        
                        ���;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     >@        ������������������������       �                     5@                                   ;@���!pc�?             &@                                    @      �?             @                                   �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @               O                    @���!pc�?4            @S@              J                    �?�w�"w��?3             S@              I                 p�w@4�2%ޑ�?/            �Q@              F                    �?�'݊U�?-            �P@              E                   �R@�����D�?+            @P@              >                    �?     8�?*             P@              )                    �?j�q����?!             I@               &                   �G@��s����?             5@              %                    �?�t����?             1@                                `f�A@؇���X�?             ,@        ������������������������       �                     �?        !       "                 @�6M@$�q-�?             *@        ������������������������       �                     @        #       $                  �}S@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        '       (                   �L@      �?             @       ������������������������       �                      @        ������������������������       �                      @        *       9                    @@д>��C�?             =@       +       .                   �@@�	j*D�?             *@        ,       -                 �̌*@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        /       6                 `f�<@z�G�z�?	             $@       0       1                 ��:@      �?              @        ������������������������       �                     @        2       3                    H@z�G�z�?             @        ������������������������       �                      @        4       5                   @L@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        7       8                   �J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        :       ;                 `fFJ@      �?
             0@       ������������������������       �                     *@        <       =                    7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ?       @                    �?؇���X�?	             ,@       ������������������������       �                     "@        A       B                    �?���Q��?             @        ������������������������       �                     �?        C       D                  x�N@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        G       H                 ���[@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        K       N                    �?r�q��?             @        L       M                  "&d@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        R       S                    (@v��:ө�?b            �c@        ������������������������       �        
             0@        T       a                    �?=��T�?X            �a@        U       ^                    �?��
ц��?	             *@       V       [                    �?���Q��?             $@       W       X                    �?      �?             @        ������������������������       �                      @        Y       Z                 `��,@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        \       ]                   �7@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        _       `                   �E@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        b       �                    �?PlX=��?O            �_@       c       �                    �?(pjm���?>            �X@       d       e                    @�q�q�?<             X@        ������������������������       �                     @        f       q                    &@f.i��n�?9            �V@        g       h                    �?D�n�3�?             3@        ������������������������       �                     @        i       p                   �P@8�Z$���?	             *@       j       o                   @H@�<ݚ�?             "@       k       n                   �5@      �?              @        l       m                   �1@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        r       s                 `f&(@��M��?-            �Q@        ������������������������       �                     @        t       u                 `f�)@�t����?*             Q@        ������������������������       �                     �?        v       �                    �?:-�.A�?)            �P@       w       �                   �*@�5��
J�?             G@       x       {                    �?l��
I��?             ;@        y       z                    ;@      �?              @        ������������������������       �                      @        ������������������������       �                     @        |       }                    @@�KM�]�?
             3@       ������������������������       �                     (@        ~                          �D@����X�?             @       ������������������������       ����Q��?             @        ������������������������       �                      @        �       �                   �2@�S����?             3@        ������������������������       �                     @        �       �                    �?z�G�z�?
             .@        ������������������������       �                     @        ������������������������       �                     (@        �       �                    �?�ՙ/�?             5@        �       �                   �7@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �@@$�q-�?             *@        �       �                   �<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     @        �       �                    :@����X�?             <@        ������������������������       �                     &@        �       �                    �?��.k���?             1@        ������������������������       �                     "@        ������������������������       �                      @        �       �                    �?��i��?           �y@        �       �                 ���.@(옄��?             G@       �       �                    �?j���� �?             A@       �       �                   �=@     ��?             @@       �       �                 P��+@      �?             <@       �       �                    �?8�A�0��?             6@        ������������������������       �                     @        �       �                   �6@     ��?             0@        �       �                 �{@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �<@z�G�z�?	             $@       �       �                 ���@�����H�?             "@        ������������������������       �                     @        �       �                   @@z�G�z�?             @       �       �                   @<@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?r�q��?             @       �       �                    �?z�G�z�?             @        ������������������������       �                     @        �       �                   �<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�8��8��?             (@        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@        �       P                   @>�y@��?�            �v@       �       �                    �?2�x���?�            @v@        �       �                    �?L
�q��?&            �M@       �       �                    �?�n_Y�K�?"             J@        �       �                  s�@�q�q�?             8@        ������������������������       �                     �?        �       �                 ���@��+7��?             7@        ������������������������       �                     @        �       �                    �?�q�q�?	             2@       �       �                 `f�@      �?             0@       �       �                   �8@�q�q�?             .@        ������������������������       �                     �?        ������������������������       �����X�?             ,@        ������������������������       �                     �?        ������������������������       �                      @        �       �                   `3@ �Cc}�?             <@       �       �                   �<@$�q-�?             :@       �       �                    �?���N8�?             5@       �       �                   �:@�X�<ݺ?             2@        ������������������������       �                     @        �       �                  s�@��S�ۿ?             .@        ������������������������       �                     @        �       �                 ��(@�C��2(�?             &@       ������������������������       �؇���X�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                    >@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 03�7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �                          �?�
dW`�?�            �r@        �       �                    @.}Z*�?.            �Q@        �       �                    �?����X�?             @        ������������������������       �                      @        �       �                 ��T?@���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        �                          �?     ��?)             P@       �       �                    �?N{�T6�?!            �K@       �       �                     @�n_Y�K�?            �C@       �       �                 ���@^H���+�?            �B@        ������������������������       �                     @        �       �                    �?      �?             @@       �       �                 ��&@R�}e�.�?             :@       �       �                    K@�q�q�?             8@       �       �                    3@�㙢�c�?             7@        �       �                    0@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 `��!@؇���X�?
             5@       �       �                 `�X!@z�G�z�?             .@       �       �                   �;@؇���X�?             ,@       �       �                    :@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    ?@r�q��?             @       ������������������������       �                     @        �       �                 `f�/@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �                         �>@      �?	             0@       �                          �*@�θ�?             *@        �       �                    <@      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @                                �;@�����H�?             "@                                 3@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @              K                0�H@����?�            @l@       	      H                   �?X�;�^o�?�            �k@       
      5                  �;@Af��?�            �j@                              ��@R�L=��?9            @X@        ������������������������       �                      @              4                   �?��K��?8            �W@                             �?�@�~6�]�?2            @U@                                �:@���H��?             E@                             �1@��(\���?             D@                             ���@؇���X�?             5@                             ���@$�q-�?             *@                              ���@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @                                �8@      �?              @                               �5@؇���X�?             @                              �?$@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     3@        ������������������������       �                      @               #                @3�@�^�����?            �E@        !      "                  �4@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        $      1                   �?��Sݭg�?            �C@       %      0                @�!@V�a�� �?             =@       &      -                pf� @�z�G��?             4@       '      (                   1@      �?	             0@        ������������������������       �      �?             @        )      ,                  �3@�8��8��?             (@        *      +                ��Y @r�q��?             @       ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     @        .      /                  �7@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     "@        2      3                   0@���Q��?             $@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@        6      G                ��y @�nkK�?H            �\@       7      F                ��) @ ,U,?��?1            �T@       8      E                   �? 7���B�?0            @T@       9      :                   ?@(�5�f��?.            �S@       ������������������������       �                    �E@        ;      <                �&B@�8��8��?             B@        ������������������������       �                     1@        =      D                @3�@�S����?             3@       >      C                  �E@�q�q�?             "@       ?      B                  �A@      �?             @       @      A                P�@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @@        I      J                   @      �?              @        ������������������������       �                     @        ������������������������       �                     @        L      M                   ;@�q�q�?             @        ������������������������       �                      @        N      O                   >@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     &@        �t�bh�h*h-K ��h/��R�(KMQKK��h]�B       �|@     �o@     �b@     �b@      O@     @T@     �N@     @T@      @      N@      �?              @      N@      �?      J@      �?      ?@      �?      �?              �?      �?                      >@              5@      @       @      @      @      @      �?              �?      @                       @              @      L@      5@     �K@      5@      K@      0@      K@      *@     �J@      (@     �J@      &@     �D@      "@      1@      @      .@       @      (@       @              �?      (@      �?      @              @      �?              �?      @              @               @       @               @       @              8@      @      "@      @      �?       @      �?                       @       @       @      @      �?      @              @      �?       @               @      �?              �?       @              �?      �?              �?      �?              .@      �?      *@               @      �?       @                      �?      (@       @      "@              @       @              �?      @      �?              �?      @                      �?      �?      �?      �?                      �?              @      �?      @      �?       @               @      �?                      @      �?              �?             �U@     �Q@              0@     �U@      K@      @      @      @      @      @      @               @      @      �?              �?      @              @      �?              �?      @              �?       @               @      �?             �S@      H@     �Q@      <@      Q@      <@      @              O@      <@      &@       @              @      &@       @      @       @      @      �?       @      �?      �?              �?      �?      @                      �?      @             �I@      4@      @              H@      4@              �?      H@      3@     �A@      &@      3@       @       @      @       @                      @      1@       @      (@              @       @      @       @       @              0@      @      @              (@      @              @      (@              *@       @      �?      @      �?                      @      (@      �?      �?      �?      �?                      �?      &@              @               @      4@              &@       @      "@              "@       @             Ps@      Z@      5@      9@      4@      ,@      2@      ,@      ,@      ,@      "@      *@              @      "@      @      �?      @      �?                      @       @       @       @      �?      @              @      �?      @      �?       @      �?      �?              �?                      �?      @      �?      @      �?      @              �?      �?      �?                      �?      �?              @               @              �?      &@      �?       @               @      �?                      "@      r@     �S@     Pq@     �S@     �C@      4@      @@      4@      @      1@      �?              @      1@              @      @      (@      @      $@      @      $@      �?              @      $@      �?                       @      9@      @      8@       @      4@      �?      1@      �?      @              ,@      �?      @              $@      �?      @      �?      @              @              @      �?              �?      @              �?      �?              �?      �?              @             �m@     �M@      F@      ;@       @      @               @       @      @       @                      @      E@      6@      A@      5@      8@      .@      8@      *@              @      8@       @      3@      @      3@      @      3@      @      �?      �?      �?                      �?      2@      @      (@      @      (@       @      @       @      @                       @       @                      �?      @                      �?               @      @      �?      @              �?      �?      �?                      �?               @      $@      @      $@      @      @      @              @      @              @                      @       @      �?      @      �?      @                      �?      @             @h@      @@      h@      <@     `g@      9@     @S@      4@               @     @S@      2@     �P@      2@     �B@      @     �B@      @      2@      @      (@      �?      @      �?      @                      �?      @              @       @      @      �?      �?      �?      �?                      �?      @                      �?      3@                       @      >@      *@      �?      @              @      �?              =@      $@      7@      @      ,@      @      (@      @      �?      @      &@      �?      @      �?      �?      �?      @              @               @       @       @                       @      "@              @      @              @      @              $@             �[@      @     �S@      @     �S@      @      S@      @     �E@             �@@      @      1@              0@      @      @      @      @      @       @       @              �?       @      �?      �?      �?      @              $@               @                       @      @@              @      @              @      @               @      @               @       @       @       @      �?              �?      &@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJf��'hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM;huh*h-K ��h/��R�(KM;��h|�B�N         f                    �?�}���?�           @�@               ]                   �?@AB����?�            `o@              "                   �2@X�Ú��?q             f@               	                     @��B����?!             J@                                   �?�	j*D�?             *@        ������������������������       �                     �?                                ���`@�q�q�?             (@       ������������������������       �                      @        ������������������������       �                     @        
                           @�e����?            �C@                                   @�	j*D�?
             *@                                  �?���|���?	             &@        ������������������������       �                     @                                P��%@և���X�?             @        ������������������������       �                      @                                    @���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @                                   (@R�}e�.�?             :@        ������������������������       �                      @                                   +@b�2�tk�?             2@        ������������������������       �                     �?                                   �?ҳ�wY;�?
             1@                               �?@����X�?             ,@        ������������������������       �                      @                                �K(@r�q��?             (@                                x&�!@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @                !                 ��'@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        #       *                    �?`�Q��?P            @_@        $       %                    �?�IєX�?             1@        ������������������������       �                      @        &       '                     @�����H�?             "@       ������������������������       �                     @        (       )                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        +       >                     @*O���?B             [@        ,       7                    �?ףp=
�?             I@       -       .                     �?\-��p�?             =@        ������������������������       �                     "@        /       6                   �7@z�G�z�?             4@       0       1                 ��Y)@���|���?             &@        ������������������������       �                     @        2       5                    �?�q�q�?             @       3       4                    :@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     "@        8       9                   �8@���N8�?             5@       ������������������������       �                     &@        :       ;                    �?ףp=
�?             $@        ������������������������       �                     @        <       =                 ���V@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ?       \                 ��Y1@�f7�z�?'             M@       @       I                    :@�`���?            �H@        A       H                    �?z�G�z�?
             .@       B       C                    �?؇���X�?	             ,@        ������������������������       �                     �?        D       G                   �6@8�Z$���?             *@       E       F                  P @�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        J       U                   �<@h+�v:�?             A@       K       T                 ��.#@l��
I��?             ;@       L       S                    �?D�n�3�?             3@       M       R                 �̌@b�2�tk�?             2@       N       O                  s�@������?	             .@        ������������������������       �                      @        P       Q                 �&B@�	j*D�?             *@       ������������������������       ����|���?             &@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        V       [                    �?����X�?             @       W       Z                   �>@���Q��?             @       X       Y                 @3#%@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        ^       _                     @�?�|�?,            �R@       ������������������������       �        (            �P@        `       c                    �?����X�?             @        a       b                    I@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        d       e                   @D@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        g       �                 `ff/@d�!��?1           �|@       h       }                    �?���H��?�            `r@        i       t                   @@R���Q�?             D@       j       k                 03S@ܷ��?��?             =@        ������������������������       �                     @        l       o                 ���@H%u��?             9@        m       n                   �7@r�q��?             (@        ������������������������       �                      @        ������������������������       �                     $@        p       s                   @<@$�q-�?	             *@       q       r                    9@�����H�?             "@        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                     @        u       x                     @���!pc�?             &@        v       w                 `��,@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        y       z                   �<@�q�q�?             @        ������������������������       �                     @        {       |                    ?@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ~                            �?�Z�)��?�            �o@        ������������������������       �                     @        �       �                   �;@��f�R@�?�            @o@        �       �                    �?��k=.��?:            �W@       �       �                    �?��3E��?9            @W@       �       �                    �?R�(CW�?4            �T@        ������������������������       �                      @        �       �                   �:@�Q��k�?3             T@       �       �                     @@�j;��?/            �Q@        �       �                    5@�t����?             1@        �       �                    &@      �?              @        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     "@        �       �                   �3@�>����?#             K@        �       �                   �2@؇���X�?             5@        �       �                 ��Y @�8��8��?             (@        �       �                 pf�@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@        �       �                 �?�@�<ݚ�?             "@        ������������������������       �                     @        �       �                 `�8"@���Q��?             @        ������������������������       ��q�q�?             @        ������������������������       �                      @        �       �                 ���@Pa�	�?            �@@        �       �                   �8@r�q��?             @       �       �                 �&b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     ;@        �       �                     @�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        �       �                 ��@���|���?             &@       ������������������������       �                     @        �       �                 �&B@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?��)�G��?e            �c@       �       �                   �<@@�+9\J�?a            �b@        ������������������������       �        %             L@        �       �                 ���@�W�{�5�?<            �W@        ������������������������       �                     1@        �       �                    �?��|��?1            �S@        �       �                   `A@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 @3�@؇���X�?-            �Q@        �       �                 �?�@     ��?             0@       �       �                   @@@ףp=
�?             $@        �       �                   �@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �D@�q�q�?             @       �       �                   �?@      �?             @        ������������������������       �                     �?        �       �                   �A@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                      @        �       �                   �"@h�WH��?              K@        ������������������������       �                     8@        �       �                   �=@r�q��?             >@        ������������������������       �                     �?        �       �                     @\-��p�?             =@       �       �                   �*@�J�4�?             9@       �       �                 `fF)@"pc�
�?             6@        �       �                 `f�&@      �?              @       �       �                   �H@؇���X�?             @       ������������������������       �                     @        �       �                   �P@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    C@d}h���?             ,@       ������������������������       �                     "@        ������������������������       ����Q��?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?h��T���?v            �d@        �       �                     �?���|���?            �@@       �       �                 @��v@r�q��?             8@       �       �                   �1@�ՙ/�?             5@        ������������������������       �                      @        �       �                 @�pX@�����?             3@       �       �                    �?�eP*L��?
             &@       �       �                 0C=@      �?	             $@        ������������������������       �                      @        �       �                  �}S@      �?              @       �       �                    �?z�G�z�?             @       �       �                 `f�B@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                 ���@@�����H�?             "@       ������������������������       �                     @        �       �                 pV�C@      �?             @       �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       $                    @.��<�?]            �`@       �                       ��YD@d�� z�?:            @T@       �                          �?�n_Y�K�?$             J@       �                          �?�"U����?#            �I@       �       �                 `fF<@b�2�tk�?             B@       �       �                   �B@r�q��?             2@        �       �                 ��$:@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                   �G@$�q-�?	             *@        ������������������������       �                     @        �       �                 `fF:@؇���X�?             @        ������������������������       �                     �?        �       �                    J@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �                          �;@b�2�tk�?
             2@        ������������������������       �                      @                                �Q@     ��?	             0@                               �J@      �?             ,@                               �H@���|���?             &@             	                �TaA@      �?              @                               �B@      �?             @                               �>@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        
                        @B@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @                                 �?�q�q�?             .@        ������������������������       �                     @                                 �?      �?             $@                                1@X�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?              #                    �?ܷ��?��?             =@                                �? �Cc}�?             <@                             03�U@HP�s��?             9@       ������������������������       �                     6@                                 �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?                                 �;@�q�q�?             @        ������������������������       �                     �?        !      "                   I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        %      0                   $@ {��e�?#            �J@        &      '                ���8@��.k���?             1@        ������������������������       �                     @        (      )                   �?ףp=
�?	             $@        ������������������������       �                     @        *      /                   @؇���X�?             @       +      .                ���A@z�G�z�?             @       ,      -                   @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        1      6                   �?�8��8��?             B@        2      5                   �?�<ݚ�?             "@       3      4                �T�C@����X�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        7      :                03�7@ 7���B�?             ;@        8      9                   �?�C��2(�?	             &@        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �        	             0@        �t�b�@     h�h*h-K ��h/��R�(KM;KK��h]�B�       |@     pp@     @Q@     �f@     �P@     �[@      ;@      9@      @      "@              �?      @       @               @      @              7@      0@      @      "@      @      @              @      @      @       @               @      @              @       @                       @      3@      @       @              &@      @              �?      &@      @      $@      @               @      $@       @      @       @      @                       @      @              �?       @               @      �?              D@     @U@      �?      0@               @      �?       @              @      �?      �?      �?                      �?     �C@     @Q@      @     �F@      @      9@              "@      @      0@      @      @              @      @       @       @       @       @                       @       @                      "@      �?      4@              &@      �?      "@              @      �?      @              @      �?              A@      8@      9@      8@      (@      @      (@       @      �?              &@       @      @       @               @      @              @                      �?      *@      5@       @      3@       @      &@      @      &@      @      &@               @      @      "@      @      @               @      @              �?                       @      @       @      @       @      @      �?      @                      �?              �?       @              "@               @      R@             �P@       @      @      �?      @      �?                      @      �?       @               @      �?             �w@     @T@     0p@     �A@      A@      @      :@      @      @              6@      @      $@       @               @      $@              (@      �?       @      �?      �?              @      �?      @               @      @      @      �?              �?      @              @       @      @              �?       @               @      �?              l@      =@      @             �k@      =@      S@      2@      S@      1@     @Q@      *@       @             �P@      *@     @P@      @      .@       @      @       @       @       @      @              "@              I@      @      2@      @      &@      �?       @      �?       @                      �?      "@              @       @      @              @       @      �?       @       @              @@      �?      @      �?      �?      �?      �?                      �?      @              ;@               @      @       @                      @      @      @      @               @      @              @       @                      �?      b@      &@     �a@      &@      L@              U@      &@      1@             �P@      &@      @      �?              �?      @              N@      $@      &@      @      "@      �?      �?      �?              �?      �?               @               @      @       @       @              �?       @      �?      �?              �?      �?               @     �H@      @      8@              9@      @              �?      9@      @      5@      @      2@      @      @      �?      @      �?      @              @      �?              �?      @              �?              &@      @      "@               @      @      @              @              @             @^@      G@      5@      (@      *@      &@      *@       @               @      *@      @      @      @      @      @       @              @      @      �?      @      �?       @               @      �?                       @       @      �?       @                      �?              �?       @                      @       @      �?      @              @      �?      �?      �?              �?      �?               @              Y@      A@      M@      7@      @@      4@      @@      3@      6@      ,@      .@      @      @       @      @                       @      (@      �?      @              @      �?      �?              @      �?              �?      @              @      &@               @      @      "@      @      @      @      @      @      @      @      �?       @      �?              �?       @              �?              �?      @              @      �?                      @      @                       @      $@      @      @              @      @      @      @              @      @              �?                      �?      :@      @      9@      @      7@       @      6@              �?       @               @      �?               @      �?      �?              �?      �?              �?      �?              �?              E@      &@      "@       @              @      "@      �?      @              @      �?      @      �?       @      �?              �?       @               @               @             �@@      @      @       @      @       @      @                       @       @              :@      �?      $@      �?              �?      $@              0@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJy"rhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM	huh*h-K ��h/��R�(KM	��h|�B@B         �                    �?�?a/���?�           @�@              �                    �?����,�?]           @�@              *                    �?���(��?           0z@                                  �5@B�����?F             Z@                                   �?
;&����?             7@                                   0@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        	                        @�"@����X�?
             ,@        
                          �4@      �?              @                               P��@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @                                    @�Zl�i��?7            @T@                                  �?p���?!             I@                                  �G@P���Q�?
             4@       ������������������������       �        	             3@        ������������������������       �                     �?        ������������������������       �                     >@               !                  ��@��a�n`�?             ?@                                  @B@R���Q�?             4@                               ���@�KM�]�?             3@                                �&�@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                  �9@�IєX�?
             1@                                  �7@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     *@        ������������������������       �                     �?        "       )                   �>@���|���?	             &@       #       $                   �8@      �?              @        ������������������������       �                     �?        %       &                   �;@և���X�?             @        ������������������������       �                      @        '       (                 @3#%@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        +       @                     �?bۘ�W^�?�            �s@        ,       ;                   �J@����3��?             J@       -       2                    �?��
P��?            �A@        .       /                 �ܵ<@      �?             $@        ������������������������       �                      @        0       1                   �A@      �?              @       ������������������������       �                     @        ������������������������       �                     @        3       :                   �>@�q�����?             9@       4       5                 ��I/@�q�q�?             2@        ������������������������       �                     @        6       9                 `fF<@$�q-�?             *@       7       8                   �A@      �?              @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        <       ?                    R@�t����?	             1@       =       >                   �@@      �?             0@       ������������������������       �                     .@        ������������������������       �                     �?        ������������������������       �                     �?        A       T                    �?����[�?�            pp@        B       I                    ;@z�G�z�?             >@        C       D                    5@      �?             @        ������������������������       �                      @        E       H                 xF*@      �?             @       F       G                 ���@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        J       Q                 pf�&@      �?             8@       K       P                    =@P���Q�?             4@       L       M                 ���@�8��8��?             (@        ������������������������       �                     @        N       O                   @@�����H�?             "@       ������������������������       �؇���X�?             @        ������������������������       �                      @        ������������������������       �                      @        R       S                 �R,@      �?             @        ������������������������       �                      @        ������������������������       �                      @        U       �                   �C@h�{��`�?�             m@       V       �                 0��D@8���|�?z            �h@       W       `                     @HKS�l�?u            �f@        X       [                    5@�˹�m��?             C@        Y       Z                   �2@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        \       ]                   �@@h�����?             <@       ������������������������       �                     4@        ^       _                   @A@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        a       �                   @C@������?^             b@       b       k                    �?���2���?\            �a@        c       d                   �:@�8��8��?             8@        ������������������������       �                     @        e       f                  s�@�t����?             1@        ������������������������       �                     @        g       j                 ��(@8�Z$���?             *@       h       i                    >@�<ݚ�?             "@       ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     @        l       q                 ��@,Z0R�?N             ]@        m       p                   �>@�q�q�?             @        n       o                 `f�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        r       �                 ���!@�o�s(��?J            �[@       s       x                 �?�@����\�?>            �V@       t       w                   �;@�&=�w��?"            �J@        u       v                    :@ףp=
�?             4@       ������������������������       �                     2@        ������������������������       �                      @        ������������������������       �                    �@@        y       �                 ��) @$G$n��?            �B@       z       {                 @3�@�����H�?             ;@        ������������������������       �r�q��?             @        |                          �3@�����?             5@        }       ~                   �1@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     2@        �       �                   �7@z�G�z�?             $@        ������������������������       �                     @        �       �                    >@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     4@        �       �                 ��	0@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    >@�	j*D�?             *@       �       �                    ;@X�<ݚ�?             "@        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                     @        �       �                   �N@�?�|�?            �B@       ������������������������       �                     A@        �       �                 hfF"@�q�q�?             @        ������������������������       �                     �?        �       �                   �P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?���)z�?R            �`@        �       �                    6@^l��[B�?$             M@        �       �                  	8@�q�q�?             (@       ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�q��/��?             G@       �       �                 pF�-@���H��?             E@        ������������������������       �                     @        �       �                     �?�7��?            �C@       ������������������������       �                     6@        �       �                     @�t����?             1@        �       �                    �?r�q��?             @        ������������������������       �                     �?        �       �                    <@z�G�z�?             @        �       �                   �7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�C��2(�?             &@        ������������������������       �                     @        �       �                 03�1@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�7�QJW�?.            �R@       �       �                    -@F�4�Dj�?&            �M@        ������������������������       �                     @        �       �                    �?X�;�^o�?%            �K@        �       �                     �?z�G�z�?             $@       �       �                   �5@���Q��?             @        ������������������������       �                     �?        �       �                 ���S@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �9@�����H�?            �F@        �       �                     @�θ�?             *@        ������������������������       �                     @        �       �                    3@�z�G��?             $@        ������������������������       �                     @        �       �                 pf(@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �>@      �?             @@        ������������������������       �                     1@        �       �                 03�U@�r����?             .@       �       �                 ��9L@@4և���?
             ,@       ������������������������       �                     &@        �       �                 03�P@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                 ���[@      �?             0@       ������������������������       �                     ,@        ������������������������       �                      @        �       �                     @R�����?k             d@       �       �                    @��C"�b�?6            �T@       �       �                    �?ڤ���?5            @T@       �       �                    �?0G���ջ?"             J@       ������������������������       �                     :@        �       �                     �?ȵHPS!�?             :@        �       �                     @���!pc�?             &@        ������������������������       �                      @        �       �                    �?�����H�?             "@       �       �                 ���`@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     .@        �       �                    �?�f7�z�?             =@        �       �                    �?      �?              @        �       �                    6@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                     �?�G��l��?             5@        �       �                     @�q�q�?             "@       �       �                   @P@      �?              @       �       �                    �?؇���X�?             @       �       �                   @K@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�q�q�?	             (@       �       �                    :@�eP*L��?             &@        ������������������������       �                     @        �       �                    $@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �                       `v�6@����[��?5            �S@       �       �                    �?4�B��?            �B@       �       �                    @"pc�
�?             6@       �       �                 ���.@ףp=
�?             4@        �       �                    �?      �?              @        ������������������������       �                     �?        �       �                   �;@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                      @        �       �                    �?��S���?             .@        ������������������������       �                     �?                                  �?և���X�?
             ,@        ������������������������       �                     @                                �1@�eP*L��?             &@                                �?؇���X�?             @                                 @r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �D@        �t�bh�h*h-K ��h/��R�(KM	KK��h]�B�        {@     �q@     `v@     @h@     �q@      a@      3@     @U@      &@      (@      @       @               @      @              @      $@      @      @      @       @               @      @                       @              @       @     @R@      �?     �H@      �?      3@              3@      �?                      >@      @      8@      @      1@       @      1@      �?      �?              �?      �?              �?      0@      �?      @              @      �?                      *@      �?              @      @      @      @      �?              @      @               @      @       @      @                       @              @     �p@     �I@     �@@      3@      2@      1@      @      @       @              @      @              @      @              *@      (@      @      (@      @              �?      (@      �?      @      �?       @              @              @      @              .@       @      .@      �?      .@                      �?              �?     �l@      @@      8@      @      @      @       @              �?      @      �?      �?              �?      �?                       @      5@      @      3@      �?      &@      �?      @               @      �?      @      �?       @               @               @       @               @       @             �i@      :@     `e@      9@     �d@      0@     �A@      @       @       @       @                       @      ;@      �?      4@              @      �?              �?      @             �`@      *@      `@      &@      6@       @      @              .@       @      @              &@       @      @       @      @       @      @              @             �Z@      "@      @       @      �?       @      �?                       @      @             �Y@      @     �T@      @     �I@       @      2@       @      2@                       @     �@@              @@      @      8@      @      @      �?      3@       @      �?       @      �?      �?              �?      2@               @       @      @              @       @               @      @              4@              @       @               @      @              @      "@      @      @              �?      @      @              @      B@      �?      A@               @      �?      �?              �?      �?              �?      �?             �R@      M@      *@     �F@       @      @       @                      @      @     �D@      @     �B@      @               @     �B@              6@       @      .@      �?      @              �?      �?      @      �?      �?      �?                      �?              @      �?      $@              @      �?      @              @      �?                      @      O@      *@      H@      &@              @      H@      @       @       @      @       @      �?               @       @               @       @              @              D@      @      $@      @      @              @      @      @              �?      @              @      �?              >@       @      1@              *@       @      *@      �?      &@               @      �?              �?       @                      �?      ,@       @      ,@                       @     �R@     �U@      5@     �N@      4@     �N@      @     �H@              :@      @      7@      @       @       @              �?       @      �?      @              @      �?                      @              .@      1@      (@      @      �?       @      �?              �?       @              @              $@      &@      @      @       @      @      �?      @      �?      @      �?                      @              @      �?              �?              @      @      @      @              @      @       @               @      @              �?              �?             �J@      9@      (@      9@      @      2@       @      2@       @      @      �?              �?      @              @      �?                      (@       @               @      @              �?       @      @      @              @      @      �?      @      �?      @              @      �?                      �?      @             �D@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�A�'hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM+huh*h-K ��h/��R�(KM+��h|�B�J         f                    �?<��z��?�           @�@               a                    @T�MB��?�            pp@              `                    @��)�?�            �m@                                  �?<��u�?�            �l@                                  �1@��|��?4            �S@        ������������������������       �        	             .@                                03�-@d�;lr�?+            �O@               	                     @      �?             8@        ������������������������       �                     @        
                           4@�G�z��?             4@        ������������������������       �                     @                                   9@     ��?             0@        ������������������������       �                      @                                   �?X�Cc�?
             ,@                                H�%@      �?             @        ������������������������       �                     �?        ������������������������       �                     @                                 ��@z�G�z�?             $@        ������������������������       �                     �?                                pF @�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?                                ��A@�7��?            �C@                                   �?      �?             0@                                `v7<@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     7@               3                     @      �?a             c@              .                 03�a@�nkK�?=             W@               !                     �?�Ń��̧?6             U@        ������������������������       �                     @@        "       -                   �;@ ��WV�?!             J@        #       ,                    �?���}<S�?             7@        $       )                    �?����X�?             @       %       &                   �'@      �?             @        ������������������������       �                     �?        '       (                   �3@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        *       +                   �9@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     0@        ������������������������       �                     =@        /       0                    �?      �?              @       ������������������������       �                     @        1       2                 Ъ�c@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        4       Q                    �?*;L]n�?$             N@       5       F                    �?Z�K�D��?            �G@       6       E                    A@��
ц��?             :@       7       <                   �5@���Q��?             4@        8       9                    3@؇���X�?             @        ������������������������       �                     @        :       ;                  P @      �?             @        ������������������������       �                     @        ������������������������       �                     �?        =       >                 pf�@��
ц��?
             *@        ������������������������       �                      @        ?       @                 �?�@���|���?             &@        ������������������������       �                     @        A       B                 `��!@և���X�?             @        ������������������������       �                     @        C       D                   P&@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        G       P                    �?���N8�?
             5@       H       O                   �=@�E��ӭ�?	             2@       I       J                 �̬)@�n_Y�K�?             *@        ������������������������       �                     @        K       L                 @3�/@r�q��?             @        ������������������������       �                     �?        M       N                    ;@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        R       [                    �?�	j*D�?
             *@       S       Z                 03S1@z�G�z�?             $@       T       Y                   �;@����X�?             @       U       X                    $@r�q��?             @       V       W                 P��%@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        \       _                    �?�q�q�?             @       ]       ^                 (C�1@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        b       c                 ��	5@ȵHPS!�?             :@        ������������������������       �                      @        d       e                      @ �q�q�?             8@        ������������������������       �                     �?        ������������������������       �        
             7@        g       p                    @Ԛ��]m�?           |@        h       i                 @3�4@�t����?             1@        ������������������������       �                     "@        j       k                    @      �?              @        ������������������������       �                     @        l       m                      @���Q��?             @        ������������������������       �                     �?        n       o                 ��T?@      �?             @        ������������������������       �                      @        ������������������������       �                      @        q       �                     �?�_p�<�?            {@        r       �                   �C@      �?8             U@       s       �                    �?�X���?              F@       t       �                    �?�4F����?            �D@        u       v                 ��>@X�Cc�?             ,@        ������������������������       �                     @        w       x                   �A@      �?             $@        ������������������������       �                      @        y       ~                    �?      �?              @       z       {                    @@      �?             @        ������������������������       �                      @        |       }                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               �                   �:@      �?             @       ������������������������       �                      @        ������������������������       �                      @        �       �                    A@l��
I��?             ;@       �       �                   �<@�GN�z�?             6@       �       �                    7@     ��?
             0@        ������������������������       �                     �?        �       �                 �̌*@�q�q�?	             .@        ������������������������       �                     @        �       �                   �;@      �?             $@        ������������������������       �                     �?        �       �                 `f�D@X�<ݚ�?             "@       �       �                   �@@�q�q�?             @       �       �                   �>@���Q��?             @       �       �                 `f�<@      �?             @       ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 ��HJ@���Q��?             @        ������������������������       �                      @        �       �                 03U@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ��^@R���Q�?             D@       �       �                    �?�?�'�@�?             C@       �       �                   �Q@��� ��?             ?@       �       �                    �?ףp=
�?             >@        �       �                   �H@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 `f�;@$�q-�?             :@        �       �                 �̌*@      �?              @        ������������������������       �                     �?        �       �                   �K@����X�?             @       �       �                    H@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     2@        ������������������������       �                     �?        �       �                 ���S@؇���X�?             @        ������������������������       �                     @        �       �                    �?      �?             @       �       �                 `��W@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                 `f�h@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �                         @@@�:���?�            �u@       �                       �T�I@vsSj��?�            �m@       �                         �3@�Fc��?�            �k@       �                         �?@ޗQ�~�?�            �i@       �       �                    +@H;T*St�?}            �h@        �       �                   X1@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�8��8��?z             h@        �       �                   �1@z�G�z�?            �A@        ������������������������       �                     @        �       �                    ;@��a�n`�?             ?@        �       �                 ���0@�	j*D�?             *@       �       �                 �{@"pc�
�?             &@        ������������������������       �                     @        �       �                    �?����X�?             @       �       �                    5@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                 ��%@r�q��?             2@       �       �                   @@�t����?
             1@       �       �                   @<@"pc�
�?             &@       �       �                 ���@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �                          �?���.n�?h            �c@       �       �                    �?�<_���?]             a@        �       �                   �<@�KM�]�?             3@       �       �                  ��@      �?             0@        ������������������������       �                      @        �       �                   @'@      �?              @       ������������������������       �r�q��?             @        ������������������������       �                      @        �       �                    >@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �<@_k,D	�?P            �]@       �       �                 ��@����?H            �Z@        �       �                     @z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �;@��'cy�?D            @Y@       �       �                     @@	tbA@�?-            @Q@        ������������������������       �        	             ,@        �       �                 @3�@ �Jj�G�?$            �K@       ������������������������       �                     <@        �       �                   �3@ 7���B�?             ;@        �       �                 ��Y @ףp=
�?             $@        �       �                   �1@      �?             @        ������������������������       �                      @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �        	             1@        �       �                  sW@     ��?             @@        �       �                 ��@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ��) @��S�ۿ?             >@       ������������������������       �                     6@        �       �                     @      �?              @        ������������������������       �                     �?        �       �                 �̜!@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                     @�q�q�?             (@        ������������������������       �                     @        �                       ���"@X�<ݚ�?             "@       �                       @3�@r�q��?             @                                 �>@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                                �9@      �?             4@              	                   7@      �?             $@                                �4@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        
                      (3�)@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     $@                                 �?      �?              @                             �?�@r�q��?             @                                �@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     3@                              p�O@և���X�?             ,@                                 >@      �?              @       ������������������������       ����Q��?             @        ������������������������       �                     @        ������������������������       �                     @                              ��)#@�?�|�?>            �[@       ������������������������       �        !             M@                                 �? �h�7W�?            �J@        ������������������������       �                      @              *                   �?�IєX�?            �I@              '                  @N@��p\�?            �D@       !      &                  @A@������?             B@        "      %                   �?؇���X�?             @       #      $                `fF)@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     =@        (      )                  �P@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     $@        �t�bh�h*h-K ��h/��R�(KM+KK��h]�B�       p|@     p@     �S@      g@      L@     �f@     �H@     �f@      &@     �P@              .@      &@      J@      "@      .@              @      "@      &@      @              @      &@               @      @      "@      @      �?              �?      @               @       @      �?              �?       @               @      �?               @     �B@       @      ,@       @      @              @       @                      "@              7@      C@     �\@      @      V@       @     �T@              @@       @      I@       @      5@       @      @      �?      @              �?      �?       @      �?      �?              �?      �?       @               @      �?                      0@              =@       @      @              @       @      �?       @                      �?      A@      :@      >@      1@      ,@      (@       @      (@      �?      @              @      �?      @              @      �?              @      @               @      @      @      @              @      @              @      @      �?      @                      �?      @              0@      @      *@      @       @      @      @              �?      @              �?      �?      @      �?                      @      @              @              @      "@       @       @       @      @      �?      @      �?       @      �?                       @              @      �?                      @       @      �?      �?      �?              �?      �?              �?              @              7@      @               @      7@      �?              �?      7@             �w@     @R@      @      (@              "@      @      @      @               @      @              �?       @       @       @                       @     0w@     �N@     �O@      5@      =@      .@      <@      *@      "@      @      @              @      @               @      @      @      @      �?       @              �?      �?      �?                      �?       @       @               @       @              3@       @      1@      @      &@      @      �?              $@      @      @              @      @              �?      @      @       @      @       @      @      �?      @      �?      �?               @      �?                      �?      @              @               @      @               @       @      �?       @                      �?      �?       @      �?                       @      A@      @     �@@      @      ;@      @      ;@      @      @      �?              �?      @              8@       @      @       @      �?              @       @      �?       @      �?      �?              �?      @              2@                      �?      @      �?      @              @      �?      �?      �?              �?      �?               @              �?      �?              �?      �?             @s@      D@      i@     �B@      h@      ?@     �e@      ?@     @e@      :@      �?      @              @      �?              e@      7@      <@      @      @              8@      @      "@      @      "@       @      @              @       @      @       @               @      @               @                       @      .@      @      .@       @      "@       @      @       @       @              @       @       @              @                      �?     �a@      0@     �_@      &@      1@       @      .@      �?       @              @      �?      @      �?       @               @      �?              �?       @             @[@      "@     @Y@      @      @      �?      @                      �?     @X@      @      Q@      �?      ,@              K@      �?      <@              :@      �?      "@      �?      @      �?       @              �?      �?      @              1@              =@      @      �?      �?      �?                      �?      <@       @      6@              @       @      �?              @       @               @      @               @      @      @              @      @      @      �?       @      �?       @                      �?      @                      @      .@      @      @      @      @      �?              �?      @               @      @              @       @              $@              @      @      �?      @      �?       @               @      �?                      @       @              3@               @      @       @      @       @      @              @      @              [@      @      M@              I@      @       @              H@      @      C@      @     �A@      �?      @      �?       @      �?      �?              �?      �?      @              =@              @       @               @      @              $@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ���hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM+huh*h-K ��h/��R�(KM+��h|�B�J                             @T�����?�           @�@               	                   p<@p9W��S�?             C@                                   �?�IєX�?             1@        ������������������������       �                     @                                �̌5@�C��2(�?             &@                                ���3@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        
                            @�G��l��?             5@                                   �?"pc�
�?             &@                                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @                                   �?z�G�z�?             $@        ������������������������       �                     @                                pf�C@����X�?             @                                  �?      �?             @                                   @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                ��T?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @               j                    �?�oMo��?�           �@               5                     �?ܐ҆��?s            @g@               4                    �?�'�`d�?*            �P@              '                 ��L@@p�v>��?            �G@               "                    �?�z�G��?             $@                !                 `v7<@      �?             @        ������������������������       �                      @        ������������������������       �                      @        #       &                   @@@r�q��?             @       $       %                 �ܵ<@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        (       -                  "�`@��G���?            �B@       )       ,                 �UP@HP�s��?             9@        *       +                  ��M@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        	             .@        .       3                 �̾w@�q�q�?	             (@       /       0                 `fpk@����X�?             @        ������������������������       �                      @        1       2                   �@@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     3@        6       i                    @��Q��?I             ^@       7       R                    �?L
�q��?H            �]@        8       O                    �?      �?             F@       9       @                    �?:ɨ��?            �@@        :       ?                   �1@      �?              @       ;       <                    0@z�G�z�?             @        ������������������������       �                      @        =       >                  Su*@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        A       B                   �2@�+e�X�?             9@        ������������������������       �                      @        C       D                   �5@��+7��?             7@        ������������������������       �                     �?        E       N                    �?�GN�z�?             6@       F       G                    9@��s����?
             5@        ������������������������       �                     @        H       M                    =@������?	             1@       I       L                 pF @      �?             0@       J       K                 ���@$�q-�?             *@        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        P       Q                 pF�-@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        S       h                    �?�����?-            �R@       T       Y                    5@ ����?*            @P@        U       V                    /@      �?              @        ������������������������       �                     �?        W       X                 �Y�@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        Z       [                    �?�}�+r��?%            �L@       ������������������������       �                     >@        \       ]                     @�����H�?             ;@        ������������������������       �                      @        ^       g                    �?H%u��?             9@       _       f                 ��(@؇���X�?             5@       `       a                  s�@z�G�z�?	             .@        ������������������������       �                     @        b       c                   �<@      �?             (@       ������������������������       �      �?              @        d       e                   �H@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                      @        k       (                   @>��/�?=           �~@       l       '                   @����V��?2           P}@       m       �                     @��J`��?+           �|@        n       �                 ��gS@4�����?�            �h@       o       �                   �K@�q�q�?w             e@       p       q                    @��&T)��?n            �b@        ������������������������       �                      @        r       }                    �?��!�^��?h            �a@        s       |                   �;@`'�J�?&            �I@        t       {                    6@�����H�?             2@        u       z                   �9@      �?              @       v       y                    �?؇���X�?             @       w       x                   �'@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �      �?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                    �@@        ~       �                     �?��wy���?B             W@               �                   �G@#z�i��?            �D@       �       �                    �?�������?             A@       �       �                   �<@      �?             @@        �       �                    7@      �?
             ,@        ������������������������       �                     �?        �       �                 ��yC@��
ц��?	             *@       �       �                   �;@�q�q�?             "@        ������������������������       �                     �?        �       �                   �@@      �?              @       �       �                   �>@���Q��?             @       �       �                 `f�<@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �;@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 03k:@�X�<ݺ?             2@        �       �                   �9@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             0@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �J@����X�?             @       �       �                   �H@r�q��?             @        ������������������������       �                     @        �       �                   @I@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?`�H�/��?&            �I@       �       �                    5@؇���X�?            �A@        �       �                    &@�q�q�?             @        �       �                   �1@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   �@@ܷ��?��?             =@       ������������������������       �                     .@        �       �                   �*@d}h���?
             ,@       �       �                   �'@�z�G��?             $@        ������������������������       �                      @        �       �                    C@      �?              @       ������������������������       �      �?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     0@        �       �                    �?�t����?	             1@        ������������������������       �                     �?        �       �                    (@      �?             0@        ������������������������       �                     �?        ������������������������       �                     .@        �       �                    4@д>��C�?             =@        �       �                    �?և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�C��2(�?             6@       ������������������������       �        	             *@        �       �                    �?�<ݚ�?             "@       �       �                    �?���Q��?             @       �       �                   �>@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       "                0��F@д>��C�?�            Pp@       �       �                    �?.vW��?�            `o@        �       �                   �K@���X�?$             L@       �       �                 �&@����|e�?#             K@        ������������������������       �                     @        �       �                    7@��x_F-�?!            �I@        �       �                    �?P���Q�?
             4@       �       �                    3@�C��2(�?             &@        �       �                 �y�+@z�G�z�?             @       �       �                 x&�!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     "@        �       �                    �?¦	^_�?             ?@       �       �                   @B@���N8�?             5@       �       �                 `�X!@�q�q�?             .@        ������������������������       �                     @        �       �                 03�1@X�<ݚ�?             "@       �       �                    ;@      �?              @        �       �                    9@      �?             @       �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 P��%@���Q��?             $@        ������������������������       �                     @        �       �                    �?և���X�?             @        ������������������������       �                      @        �       �                     @���Q��?             @       �       �                 03S1@      �?             @        ������������������������       �                     �?        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       !                   �?�?�<��?y            `h@       �                        ��i @H�g�}N�?q            �f@       �                         �F@:	��ʵ�?S            �`@       �                         �E@�2�KZ�?J            @^@       �                         @@@�V�i�#�?I            @]@       �                         �?@�\m����?;             Y@       �                         �>@v�9�z��?:            @X@       �                         �<@�S����?8            �W@       �                         �:@r�q��?5            �V@       �                         �9@؇���X�?              L@       �                          �?�㙢�c�?             G@       �                         �5@X�EQ]N�?            �E@       �       �                 @3�@�חF�P�?             ?@       �       �                 �1@���N8�?             5@        �       �                    4@ףp=
�?             $@       ������������������������       �                      @        �       �                  s@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     &@                                 �3@���Q��?             $@                               �1@X�<ݚ�?             "@        ������������������������       ����Q��?             @        ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                     @        ������������������������       �                     $@              	                  �;@H�V�e��?             A@        ������������������������       �                      @        
                         �?     ��?             @@                             ��) @r�q��?             >@                             �?$@ �Cc}�?             <@                              pf�@      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     6@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @                              pff@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                              �?�@�IєX�?             1@        ������������������������       �                     "@                              @3�@      �?              @                                 �?�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        	             ,@        ������������������������       �                    �G@        ������������������������       �                     *@        #      &                   >@���Q��?             $@       $      %                   ;@և���X�?             @        ������������������������       �                      @        ������������������������       �z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     &@        )      *                ���3@�}�+r��?             3@        ������������������������       �                     �?        ������������������������       �        
             2@        �t�b�      h�h*h-K ��h/��R�(KM+KK��h]�B�       0|@     Pp@      &@      ;@      �?      0@              @      �?      $@      �?      @              @      �?                      @      $@      &@       @      "@       @       @       @                       @              @       @       @      @              @       @       @       @      �?      �?      �?                      �?      �?      �?      �?                      �?      @             �{@     @m@      W@     �W@      ,@      J@      ,@     �@@      @      @       @       @               @       @              @      �?      @      �?      @                      �?       @              @      >@       @      7@       @       @               @       @                      .@      @      @      @       @       @              @       @      @                       @              @              3@     �S@      E@     �S@      D@      &@     �@@      $@      7@      @      @      �?      @               @      �?       @               @      �?              @              @      3@               @      @      1@      �?              @      1@      @      1@              @      @      *@      @      (@      �?      (@      �?                      (@      @                      �?      �?              �?      $@      �?                      $@     �P@      @      M@      @      @      @              �?      @      @      @                      @      K@      @      >@              8@      @       @              6@      @      2@      @      (@      @      @              "@      @      @      �?       @       @               @       @              @              @              "@                       @     �u@     �a@     �t@     `a@     �s@     `a@     �Y@     �W@     �X@     �Q@     �T@      Q@       @             �R@      Q@       @     �H@       @      0@       @      @      �?      @      �?      @              �?      �?      @               @      �?                      $@             �@@     @R@      3@      ;@      ,@      9@      "@      8@       @      @      @      �?              @      @      @      @              �?      @      @      @       @       @       @       @      �?              �?      �?                      @      @      �?              �?      @              1@      �?      �?      �?      �?                      �?      0@              �?      �?      �?                      �?       @      @      �?      @              @      �?       @      �?                       @      �?              G@      @      >@      @      @       @      �?       @      �?                       @      @              :@      @      .@              &@      @      @      @       @              @      @      @      @       @              @              0@              .@       @              �?      .@      �?              �?      .@              @      8@      @      @              @      @               @      4@              *@       @      @       @      @      �?      @      �?                      @      �?                      @      k@     �F@     �j@     �C@     �D@      .@     �D@      *@              @     �D@      $@      3@      �?      $@      �?      @      �?      �?      �?      �?                      �?      @              @              "@              6@      "@      0@      @      $@      @      @              @      @      @      @      @      �?      �?      �?      �?                      �?       @                      @      �?              @              @      @      @              @      @               @      @       @       @       @      �?              �?       @               @      �?              �?                       @     `e@      8@     �c@      8@     �[@      8@     @X@      8@     @X@      4@     @T@      3@     @T@      0@      T@      .@     �R@      .@      H@       @      C@       @      C@      @      :@      @      4@      �?      "@      �?       @              �?      �?      �?                      �?      &@              @      @      @      @      @       @       @       @      �?              (@                      @      $@              ;@      @               @      ;@      @      9@      @      9@      @      @      @      @                      @      6@                       @       @              @              �?      �?      �?                      �?              @      0@      �?      "@              @      �?       @      �?      �?      �?      �?              @                      @      ,@             �G@              *@              @      @      @      @               @      @      �?              @      &@              2@      �?              �?      2@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJJ��hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM9huh*h-K ��h/��R�(KM9��h|�B@N         n                     @�)�>_M�?�           @�@               #                    �?և���X�?�            �r@                                   @t�e�í�?R            �`@        ������������������������       �                     @                                    �?�Ώ��?Q            ``@                               ���a@�ӖF2��?*            �Q@                                  �?���U�?"            �L@               	                   �H@      �?             @@       ������������������������       �                     7@        
                           �?�<ݚ�?             "@                                   �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     9@                                03c@d}h���?             ,@        ������������������������       �                     @        ������������������������       �                     &@               "                    �?(;L]n�?'             N@              !                   �;@h�����?$             L@                                  �?@4և���?             <@        ������������������������       �                     @                                   �?�C��2(�?             6@                                 �6@�����H�?             "@        ������������������������       �                     @                                  �8@      �?             @                                  �?�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                    6@$�q-�?             *@        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                     <@        ������������������������       �                     @        $       %                    &@�|G7�?p            �d@        ������������������������       �                     $@        &       m                    �?�&z{�?k            �c@       '       V                     �?�S���Q�?e            �b@       (       E                   �E@�e����?4            �S@       )       4                   �>@      �?              F@        *       +                 ��$:@�z�G��?             4@        ������������������������       �                     @        ,       1                    B@      �?             0@       -       0                 �ܵ<@$�q-�?             *@        .       /                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     &@        2       3                   �C@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        5       6                  x#J@�q�q�?             8@        ������������������������       �                      @        7       8                   �8@      �?             0@        ������������������������       �                     @        9       :                    <@�q�q�?
             (@        ������������������������       �                     @        ;       <                    >@X�<ݚ�?             "@        ������������������������       �                      @        =       >                 03�P@����X�?             @        ������������������������       �                     @        ?       @                    �?      �?             @        ������������������������       �                     �?        A       B                 03U@�q�q�?             @        ������������������������       �                     �?        C       D                 ��n^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        F       G                   �G@�t����?             A@        ������������������������       �                      @        H       K                 ���=@�n_Y�K�?             :@        I       J                   �J@8�Z$���?             *@        ������������������������       �                      @        ������������������������       �                     &@        L       S                    �?�n_Y�K�?             *@       M       P                    �?      �?              @        N       O                   �K@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        Q       R                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        T       U                 03�S@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        W       j                    M@@�j;��?1            �Q@       X       ]                    4@�IєX�?/             Q@        Y       \                    �?z�G�z�?             $@       Z       [                    &@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ^       i                    �?XB���?)             M@       _       h                    =@ �#�Ѵ�?            �E@       `       g                    �?HP�s��?             9@       a       b                   �'@�8��8��?             8@        ������������������������       �                      @        c       f                   �*@      �?	             0@       d       e                   �:@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     2@        ������������������������       �                     .@        k       l                   �P@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        o       �                    �?�:���?           �y@        p       y                 ���@t�Hr;��?L            ``@        q       t                    �?      �?	             0@        r       s                   �0@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        u       v                 ��Y@$�q-�?             *@        ������������������������       �                     @        w       x                   �7@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        z       �                    �?���Q��?C            �\@        {       �                 ���.@      �?             H@       |       �                    �?H�z�G�?             D@        }       �                    �?      �?             (@       ~                           .@�q�q�?             "@        ������������������������       �                     @        �       �                 ���%@���Q��?             @        ������������������������       �                     �?        �       �                   �<@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    ?@��>4և�?             <@       �       �                    �?�G��l��?             5@       �       �                    �?�G�z��?
             4@       �       �                 H�Z&@�\��N��?	             3@       �       �                   @@j���� �?             1@       �       �                   @<@�q�q�?             (@       �       �                    5@      �?             $@        ������������������������       �                     �?        �       �                    9@X�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �և���X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?      �?              @       �       �                    �?z�G�z�?             @        �       �                   �2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?��y�:�?'            �P@        �       �                    �?���@M^�?             ?@       �       �                    �?J�8���?             =@       �       �                   �2@���Q��?             9@        ������������������������       �                     @        �       �                 pF @�G��l��?             5@       �       �                   �5@b�2�tk�?
             2@        ������������������������       �                     @        �       �                 ���@������?	             .@        ������������������������       �                     �?        �       �                 ���@d}h���?             ,@        ������������������������       �                     @        �       �                    9@�z�G��?             $@        ������������������������       �                     @        �       �                 �&B@և���X�?             @       ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                 03�7@�8��8��?             B@       �       �                   �=@ܷ��?��?             =@       �       �                   `3@r�q��?             2@       �       �                   �8@�t����?             1@        ������������������������       �                     @        �       �                 ��(@؇���X�?
             ,@       �       �                 03�@z�G�z�?             $@        ������������������������       �                      @        �       �                    �?      �?              @       ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     @        �       �                    �?������?�            �q@        �       �                 �&B@��cv�?4            @S@        �       �                 ���@ףp=
�?             $@       ������������������������       �                     @        �       �                   �7@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                 `f7@��ga�=�?.            �P@       �       �                    @��V#�?            �E@       �       �                    �?������?            �D@       �       �                    �?�d�����?             C@        �       �                   �;@R���Q�?             4@       �       �                    �?���!pc�?             &@       �       �                    3@      �?              @        �       �                 x&�!@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    -@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        �       �                    �?b�2�tk�?             2@       �       �                    ;@��
ц��?	             *@        ������������������������       �                     @        �       �                     @؇���X�?             @       �       �                   �D@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    >@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 �̌5@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    �? �q�q�?             8@        ������������������������       �                     @        �       �                    @�X�<ݺ?             2@        ������������������������       �                     "@        �       �                    @�����H�?             "@        �       �                 ��T?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @��9~��?�            `i@        �       �                 pf�C@      �?              @       ������������������������       �                     @        ������������������������       �                     @        �       8                   �?�ݜ�?�            `h@       �       1                  @@@$�{�F"�?w             e@       �       ,                ��C@\|/��j�?]            �`@       �       �                 ��@̌WZ�}�?X            �^@        �       �                    6@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       	                  �4@�^����?U            �]@        �       �                   �0@      �?             4@        �       �                 pf�@���Q��?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        �                          �2@z�G�z�?             .@        ������������������������       �                     @                                �3@�q�q�?             "@                             pf�@�q�q�?             @        ������������������������       �                     @                              `�8"@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                 �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        
      !                  �>@�)���Y�?G            �X@                             �1@t��ճC�?>             V@                              �?$@PN��T'�?             ;@                               �8@�nkK�?             7@                                 7@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     1@                                �8@      �?             @        ������������������������       �                     �?        ������������������������       �                     @                                �:@�]0��<�?/            �N@        ������������������������       �                     7@                                  �?�}�+r��?             C@                               �;@      �?             @@        ������������������������       �                     �?                                @<@�g�y��?             ?@                             ��) @�nkK�?             7@       ������������������������       �                     2@                              pf� @z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        "      +                ��I @�z�G��?	             $@       #      &                  �?@      �?              @        $      %                pff@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        '      (                  �@�q�q�?             @        ������������������������       �                     �?        )      *                �?�@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �      �?             @        ������������������������       �                      @        -      0                   >@�q�q�?             "@       .      /                   ;@և���X�?             @        ������������������������       �                     �?        ������������������������       �      �?             @        ������������������������       �                      @        2      3                  �E@@-�_ .�?            �B@       ������������������������       �                     5@        4      7                @3�@      �?             0@       5      6                   G@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     :@        �t�bh�h*h-K ��h/��R�(KM9KK��h]�B�       `{@      q@      `@     �e@      $@      _@      @              @      _@      @     �P@       @     �K@       @      >@              7@       @      @       @      �?       @                      �?              @              9@      @      &@      @                      &@       @      M@       @      K@       @      :@              @       @      4@      �?       @              @      �?      @      �?       @      �?      �?              �?              �?      �?      (@      �?                      (@              <@              @     �]@      H@              $@     �]@      C@     �[@      C@      G@      @@      6@      6@      @      ,@      @               @      ,@      �?      (@      �?      �?      �?                      �?              &@      �?       @      �?                       @      0@       @       @               @       @      @              @       @              @      @      @       @               @      @              @       @       @              �?       @      �?      �?              �?      �?              �?      �?              8@      $@       @              0@      $@      &@       @               @      &@              @       @       @      @      �?      @      �?                      @      �?       @               @      �?              @       @               @      @             @P@      @      P@      @       @       @      @       @               @      @               @              L@       @     �D@       @      7@       @      6@       @       @              ,@       @       @       @       @                       @      @              �?              2@              .@              �?       @               @      �?               @             Ps@     �Y@     �T@      H@      ,@       @       @      �?              �?       @              (@      �?      @              @      �?              �?      @             @Q@      G@      8@      8@      7@      1@      @      @      @      @              @      @       @              �?      @      �?      @                      �?      @              1@      &@      $@      &@      "@      &@      "@      $@      @      $@      @      @      @      @              �?      @      @       @              @      @       @                      @       @                      �?      �?              @              �?      @      �?      @      �?      �?      �?                      �?              @              @     �F@      6@      (@      3@      $@      3@      $@      .@              @      $@      &@      @      &@      @              @      &@      �?              @      &@              @      @      @              @      @      @      @      @              �?      @                      @       @             �@@      @      :@      @      .@      @      .@       @      @              (@       @       @       @       @              @       @      @       @       @              @                      �?      &@              @             @l@      K@     �J@      8@      �?      "@              @      �?      @              @      �?              J@      .@      =@      ,@      =@      (@      <@      $@      1@      @       @      @      @      �?      @      �?      @                      �?      @              �?       @      �?                       @      "@              &@      @      @      @      @              �?      @      �?      @              @      �?                       @      @      �?      @                      �?      �?       @      �?                       @               @      7@      �?      @              1@      �?      "@               @      �?      �?      �?      �?                      �?      @             �e@      >@      @      @              @      @             @e@      9@      b@      9@     @[@      7@     �Z@      1@       @      @       @                      @      Z@      ,@      .@      @      @       @       @              �?       @      (@      @      @              @      @      @       @      @              �?       @               @      �?               @      �?       @                      �?     @V@      "@     �T@      @      7@      @      6@      �?      @      �?      @                      �?      1@              �?      @      �?                      @     �M@       @      7@              B@       @      >@       @              �?      >@      �?      6@      �?      2@              @      �?              �?      @               @              @              @      @      @      @      �?      �?      �?                      �?      @       @              �?      @      �?      �?              @      �?       @              @      @      @      @              �?      @      @               @     �A@       @      5@              ,@       @      @       @               @      @               @              :@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�U�uhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM)huh*h-K ��h/��R�(KM)��h|�B@J         r                     @r�����?�           @�@                                   �?� �	��?�            Pt@                                03[=@����?�?Q            �`@                                   �?����˵�?#            �M@                                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @                                  �+@@3����?             K@        	       
                 `f�)@���N8�?             5@        ������������������������       �                     @                                   :@��S�ۿ?             .@        ������������������������       �z�G�z�?             @        ������������������������       �                     $@        ������������������������       �                    �@@        ������������������������       �        .             S@               K                     �?�d�����?y            �g@                                  2@uvI��?>            �X@        ������������������������       �                     @               $                    �?�x�(��?;             W@               #                   �J@�5��?             ;@                                  �?8����?             7@                                  �?������?             1@                               ���<@����X�?	             ,@        ������������������������       �                     @                                  �C@X�<ݚ�?             "@                               ���Z@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @               "                   �H@      �?             @               !                 ���X@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        %       F                    �?�	j*D�?)            @P@       &       =                    �?��N`.�?!            �K@       '       <                    R@��]�T��?            �D@       (       ;                   @J@�q�q�?            �C@       )       4                   �>@     ��?             @@       *       -                    A@և���X�?             5@        +       ,                 `fF<@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        .       /                   �E@����X�?             ,@        ������������������������       �                     @        0       1                 ��:@X�<ݚ�?             "@        ������������������������       �                      @        2       3                    H@����X�?             @       ������������������������       ����Q��?             @        ������������������������       �                      @        5       :                   �=@�C��2(�?             &@       6       9                 `f�D@r�q��?             @        7       8                   �@@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        >       ?                    <@d}h���?	             ,@        ������������������������       �                     �?        @       E                    D@8�Z$���?             *@        A       B                    >@����X�?             @        ������������������������       �                     @        C       D                   @K@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        G       J                   �B@z�G�z�?             $@        H       I                   �<@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        L       e                    �?��A��?;             W@       M       N                    !@�����H�?*            �O@        ������������������������       �                     �?        O       d                   �*@��a�n`�?)             O@       P       Q                    @�t����?            �I@        ������������������������       �                     @        R       ]                   @C@��E�B��?            �G@       S       Z                    @@ >�֕�?            �A@       T       Y                    5@h�����?             <@        U       X                    &@      �?              @        V       W                   �1@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     4@        [       \                   �'@؇���X�?             @        ������������������������       �                      @        ������������������������       �z�G�z�?             @        ^       _                   �F@�q�q�?             (@        ������������������������       �      �?             @        `       c                 `f'@      �?              @        a       b                   �P@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        
             &@        f       g                    +@V�a�� �?             =@        ������������������������       �                     @        h       i                    �? �q�q�?             8@        ������������������������       �                      @        j       q                    :@���7�?
             6@       k       l                   �<@�8��8��?             (@        ������������������������       �                     @        m       n                   �7@r�q��?             @        ������������������������       �                      @        o       p                   �@@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        s       (                   @���t�?�            0x@       t       �                 `f�%@����X�?�            0w@       u       �                 pF @�Z�LY�?�            �n@       v       �                    �?� <�+�?m            �d@       w       x                    +@H�z�'�?l             d@        ������������������������       �                      @        y       �                 03�@�@G���?k            �c@        z       {                    �?�}�+r��?             3@        ������������������������       �                     @        |       }                    :@$�q-�?	             *@       ������������������������       �                     $@        ~                        ��@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?�^�!<�?`            `a@        �       �                    �?^��>�b�?*            @P@        �       �                    �?������?             ;@        ������������������������       �                     @        �       �                 �&B@�q�q�?             5@       �       �                 ���@j���� �?	             1@        �       �                 ���@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �5@���Q��?             $@        ������������������������       �                      @        �       �                    9@      �?              @        ������������������������       �                     �?        ������������������������       �և���X�?             @        ������������������������       �                     @        �       �                    �?���y4F�?             C@       �       �                   �7@�<ݚ�?             B@        �       �                 ���@����X�?             @       �       �                 ���@r�q��?             @        ������������������������       �                     @        �       �                    5@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?ܷ��?��?             =@       �       �                   @<@8�Z$���?             *@       �       �                   �:@z�G�z�?	             $@        ������������������������       �                     �?        �       �                 ���@�<ݚ�?             "@        ������������������������       �                     @        �       �                   @@�q�q�?             @       ������������������������       ����Q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ��(@      �?
             0@       �       �                 03�@@4և���?	             ,@        ������������������������       �                     �?        �       �                   �<@$�q-�?             *@        ������������������������       �                      @        �       �                   �>@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?�MI8d�?6            �R@       �       �                 �?�@r�q��?4             R@       �       �                    �?X��Oԣ�?,             O@       �       �                   �;@�KM�]�?(            �L@        �       �                   �:@r�q��?             >@       �       �                 ���@ �Cc}�?             <@        �       �                 ���@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �? �q�q�?             8@        �       �                    2@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     4@        ������������������������       �                      @        �       �                    =@ 7���B�?             ;@       �       �                 �?$@�IєX�?             1@        �       �                 pf�@؇���X�?             @       ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     $@        ������������������������       �                     $@        �       �                   �7@z�G�z�?             @        ������������������������       �                     @        �       �                   �9@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?      �?             $@       �       �                   �:@X�<ݚ�?             "@        ������������������������       �                      @        �       �                   �D@����X�?             @       �       �                   �A@�q�q�?             @        ������������������������       �      �?             @        ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?ףp=
�?4             T@       �       �                  �#@���Lͩ�?1            �R@       �       �                   �0@@4և���?.            �Q@        �       �                 pFD!@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        �       �                    �?���7�?+            �P@       �       �                 pf!@P���Q�?'             N@        ������������������������       �                     <@        �       �                   �>@     ��?             @@       �       �                 ���!@���7�?             6@       �       �                    8@ףp=
�?             $@       ������������������������       �                     @        �       �                   �;@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        �       �                    �?z�G�z�?             $@        �       �                  SE"@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                 03$@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    $@z�G�z�?             @        ������������������������       �                      @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 pf�+@xk�2���?H            �_@        ������������������������       �                     &@        �       �                 `�X.@J�8���?B             ]@        ������������������������       �        	             .@        �                       03c4@D��ٝ�?9            @Y@        �                          �?�n_Y�K�?            �C@       �       �                 03�1@r�q��?             8@       �       �                    �?��S�ۿ?	             .@       �       �                 @3�/@�8��8��?             (@        ������������������������       �                     @        �       �                    ;@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                                  �?�q�q�?             "@        ������������������������       �                     �?                               �2@      �?              @        ������������������������       �                     @        ������������������������       �                     @              
                   �?������?	             .@              	                   �?      �?             @                               �2@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?                                 0@�����H�?             "@                              `ff/@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @                                 �?r֛w���?!             O@                                 �?��.k���?
             1@        ������������������������       �                     �?                                 >@     ��?	             0@                                ;@      �?             (@                                 �?      �?             @        ������������������������       �                      @        ������������������������       �                      @                                 �?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @              !                   @:	��ʵ�?            �F@                                 @`2U0*��?             9@                              �̌5@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     7@        "      #                ��T?@��Q��?
             4@        ������������������������       �                     @        $      %                   �?��
ц��?             *@        ������������������������       �                     @        &      '                   @�z�G��?             $@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     0@        �t�bh�h*h-K ��h/��R�(KM)KK��h]�B�       �z@      r@     �a@     �f@      @     �`@      @      L@       @      @       @                      @      �?     �J@      �?      4@              @      �?      ,@      �?      @              $@             �@@              S@     �a@      I@     �N@     �B@              @     �N@      ?@      0@      &@      0@      @      *@      @      $@      @      @              @      @      @      @              @      @               @              @              @      @      �?      @              @      �?               @                      @     �F@      4@     �B@      2@      :@      .@      :@      *@      3@      *@      "@      (@      @       @      @                       @      @      $@              @      @      @       @               @      @       @      @               @      $@      �?      @      �?       @      �?       @                      �?      @              @              @                       @      &@      @              �?      &@       @      @       @      @              �?       @      �?                       @      @               @       @      @       @      @                       @      @             �S@      *@      L@      @              �?      L@      @     �F@      @      @             �D@      @     �@@       @      ;@      �?      @      �?      @      �?      �?               @      �?      @              4@              @      �?       @              @      �?       @      @      �?      @      @      �?       @      �?              �?       @              @              &@              7@      @              @      7@      �?       @              5@      �?      &@      �?      @              @      �?       @              @      �?              �?      @              $@             �q@     �Z@     �p@     �Z@     �g@     �K@     @]@     �G@     @]@     �E@               @     @]@     �D@      2@      �?      @              (@      �?      $@               @      �?       @                      �?     �X@      D@     �B@      <@      @      4@              @      @      ,@      @      $@      �?      @      �?                      @      @      @       @              @      @              �?      @      @              @      >@       @      <@       @       @      @      �?      @              @      �?       @               @      �?              �?              :@      @      &@       @       @       @      �?              @       @      @              @       @      @       @      �?              @              .@      �?      *@      �?      �?              (@      �?       @              @      �?              �?      @               @               @              O@      (@      N@      (@     �K@      @     �I@      @      9@      @      9@      @       @       @       @                       @      7@      �?      @      �?      @                      �?      4@                       @      :@      �?      0@      �?      @      �?      @              �?      �?      $@              $@              @      �?      @              �?      �?              �?      �?              @      @      @      @       @               @      @       @      @      �?      @      �?      �?              �?      �?               @                      @      R@       @      Q@      @     @P@      @       @       @      �?       @      �?             �O@      @     �L@      @      <@              =@      @      5@      �?      "@      �?      @              @      �?              �?      @              (@               @       @      @       @               @      @              @              @              @       @               @      @              @      �?       @               @      �?              �?       @              S@     �I@              &@      S@      D@      .@             �N@      D@      .@      8@      @      4@      �?      ,@      �?      &@              @      �?      @      �?                      @              @      @      @              �?      @      @      @                      @      &@      @      @      @       @      @       @                      @      �?               @      �?      @      �?      @                      �?      @              G@      0@      "@       @              �?      "@      @      "@      @       @       @               @       @              @      �?      @                      �?              @     �B@       @      8@      �?      �?      �?      �?                      �?      7@              *@      @      @              @      @      @              @      @              @      @              0@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJW��]hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM	huh*h-K ��h/��R�(KM	��h|�B@B         L                    �?�Qc�!�?�           @�@               C                    @ڤ���?�            `n@              
                    �?�b<�J�?�            �k@                                    @ pƵHP�?             J@       ������������������������       �                    �A@                                P��+@�IєX�?
             1@        ������������������������       �                     "@               	                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     @                                    @�&�+�?k            `e@                               ���`@hl �&�?=             W@                                 �+@����ȫ�?6            �T@                                  �9@ �q�q�?             8@                                  �'@z�G�z�?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                     3@        ������������������������       �        &             M@                                   ;@z�G�z�?             $@                                   �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                ���@bf@����?.            �S@        ������������������������       �                      @               (                   �9@:%�[��?(            �Q@               !                  �#@V�a�� �?             =@                                   �?�X�<ݺ?	             2@                                  �5@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     .@        "       #                  �M$@�eP*L��?             &@        ������������������������       �                      @        $       '                    �?�q�q�?             "@       %       &                 hVE0@���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        )       6                   �<@�G��l��?             E@       *       +                    @���N8�?             5@       ������������������������       �        	             $@        ,       /                    �?�eP*L��?             &@        -       .                 03�'@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        0       1                   �*@�q�q�?             @        ������������������������       �                      @        2       3                   �.@      �?             @        ������������������������       �                     �?        4       5                    ;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        7       B                   �K@����X�?	             5@       8       =                    �?      �?             4@        9       <                   �@@���|���?             &@        :       ;                 @3#%@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        >       ?                 `f�/@�����H�?             "@        ������������������������       �                     @        @       A                   �@@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        D       E                 ��	5@��Q��?             4@        ������������������������       �                     @        F       G                      @     ��?             0@        ������������������������       �                      @        H       K                    @@4և���?
             ,@        I       J                    @�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        M       �                     �?>��O�V�?*           P}@        N       �                    �?և���X�?>            �X@       O       �                 ��^@���3E��?:            @W@       P       �                    �?\�G�2��?6            @U@       Q       �                    �?\�Uo��?1             S@       R       Y                    �?�Gi����?0            �R@        S       T                   �;@և���X�?	             ,@        ������������������������       �                     @        U       V                 ��hU@�����H�?             "@       ������������������������       �                     @        W       X                 @�pX@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        Z       q                    �?���Q��?'             N@       [       j                   �>@�û��|�?             G@       \       i                    R@      �?             A@       ]       ^                   �9@`՟�G��?             ?@        ������������������������       �                     @        _       h                   �J@�q�q�?             8@       `       g                   `G@@�0�!��?             1@       a       b                 03k:@���!pc�?             &@        ������������������������       �                     @        c       f                   @>@      �?              @       d       e                   �<@���Q��?             @        ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        k       p                   �=@�8��8��?             (@       l       o                 ��yC@r�q��?             @        m       n                   �@@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        r                           D@և���X�?
             ,@       s       ~                   �B@�eP*L��?             &@       t       }                   �@@X�<ݚ�?             "@       u       v                 `fFJ@և���X�?             @        ������������������������       �                     �?        w       |                    >@�q�q�?             @       x       {                 ���M@�q�q�?             @       y       z                    7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�����H�?             "@        ������������������������       �                     @        �       �                    �?r�q��?             @        ������������������������       �                     @        �       �                 Ј�P@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?      �?              @       �       �                    �?r�q��?             @       �       �                   �<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                 �̰f@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    *@࿖��H�?�            0w@        �       �                     @      �?             4@       �       �                    $@r�q��?             (@       ������������������������       �                      @        �       �                    '@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?�6L��?�            �u@       �       �                   �<@Tri����?�            �q@       �       �                 ���@��;M��?q            @f@        �       �                    �?���N8�?             5@        �       �                 ��Y@"pc�
�?             &@        ������������������������       �                     @        �       �                   �7@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                 �&b@�z�G��?             $@       �       �                   �:@      �?              @        �       �                   �6@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                     @�B�ǈ�?c            �c@        �       �                    �?�IєX�?             A@        ������������������������       �                      @        �       �                   �;@      �?             @@       �       �                    5@�g�y��?             ?@        �       �                   �2@�C��2(�?             &@       ������������������������       �                     "@        �       �                   �'@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        
             4@        ������������������������       �                     �?        �       �                 �T)D@@;�"�?P            �^@       �       �                   �;@�IєX�?M            �]@        �       �                    �?�8��8��?&             N@        ������������������������       �                      @        �       �                 ���!@��ϭ�*�?%             M@       �       �                 @3�@�q��/��?             G@       �       �                   �5@ �q�q�?             8@       �       �                 �1@@4և���?	             ,@        �       �                 �?$@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     $@        �       �                 pf� @"pc�
�?             6@       �       �                   �3@"pc�
�?             &@        �       �                   �1@���Q��?             @       ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �7@"pc�
�?             &@       ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                     (@        �       �                    �?���#�İ?'            �M@        ������������������������       �                     3@        �       �                 �?$@P���Q�?             D@        �       �                 pf�@r�q��?             @       ������������������������       �                     @        ������������������������       ��q�q�?             @        �       �                 ��) @г�wY;�?             A@       ������������������������       �                     5@        �       �                 pf� @$�q-�?             *@        ������������������������       �                     �?        ������������������������       �                     (@        �       �                    ;@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 0��D@�ջ����?A             Z@       �       �                    �?�DÓ ��??            @Y@        ������������������������       �                     "@        �       �                     @*
;&���?:             W@        �       �                   @A@XB���?             =@        �       �                   �@@�����H�?             "@        ������������������������       �                     @        ������������������������       �z�G�z�?             @        ������������������������       �        
             4@        �       �                   �=@Z���c��?*            �O@        �       �                    �?r�q��?             @        ������������������������       �                     �?        �       �                 �̌!@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 @3�@Ԫ2��?'            �L@       �       �                   @F@r٣����?            �@@       �       �                   �E@�	j*D�?             :@       �       �                 �?�@      �?             8@       �       �                   �@@�X�<ݺ?             2@        �       �                    �?�����H�?             "@        ������������������������       �                     @        �       �                 �&B@      �?             @        ������������������������       �                      @        �       �                   �@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        �       �                   �A@r�q��?             @       ������������������������       �z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     8@        ������������������������       �                     @        �                            @�nkK�?,            @Q@        ������������������������       �                     1@                                 �?0G���ջ?              J@                                �1@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                              �&B@`2U0*��?             I@                              ��@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                    �F@        �t�b��     h�h*h-K ��h/��R�(KM	KK��h]�B�       �{@     �p@      N@     �f@     �G@      f@      �?     �I@             �A@      �?      0@              "@      �?      @      �?                      @      G@     @_@      @     @V@      �?     @T@      �?      7@      �?      @               @      �?       @              3@              M@       @       @       @      �?              �?       @                      @     �E@      B@               @     �E@      <@      7@      @      1@      �?       @      �?       @                      �?      .@              @      @               @      @      @       @      @       @                      @      @              4@      6@      @      0@              $@      @      @      @       @      @                       @       @      @               @       @       @      �?              �?       @      �?                       @      .@      @      .@      @      @      @      @      @      @                      @      @               @      �?      @               @      �?       @                      �?              �?      *@      @              @      *@      @               @      *@      �?       @      �?       @                      �?      &@             �w@     �U@      L@      E@     �K@      C@      K@      ?@      G@      >@      F@      >@       @      @              @       @      �?      @              �?      �?              �?      �?              B@      8@      <@      2@      1@      1@      1@      ,@      @              $@      ,@      @      ,@      @       @              @      @      @      @       @      �?       @       @                      @              @      @                      @      &@      �?      @      �?      �?      �?      �?                      �?      @              @               @      @      @      @      @      @      @      @      �?               @      @       @      �?      �?      �?      �?                      �?      �?                      @       @                       @      @               @               @      �?      @              @      �?      @               @      �?              �?       @              �?      @      �?      @      �?       @      �?                       @              @               @      �?      @              @      �?             `t@     �F@      $@      $@       @      $@               @       @       @       @                       @       @             �s@     �A@     @o@      @@     `d@      .@      0@      @      "@       @      @              @       @               @      @              @      @      @      �?       @      �?       @                      �?      @                       @     `b@      $@      @@       @       @              >@       @      >@      �?      $@      �?      "@              �?      �?              �?      �?              4@                      �?     �\@       @      \@      @     �K@      @       @             �J@      @     �D@      @      7@      �?      *@      �?      @      �?      @                      �?      $@              $@              2@      @      "@       @      @       @      @      �?              �?      @              "@       @      "@                       @      (@             �L@       @      3@              C@       @      @      �?      @               @      �?     �@@      �?      5@              (@      �?              �?      (@              @      �?              �?      @             �U@      1@     �U@      ,@      "@             �S@      ,@      <@      �?       @      �?      @              @      �?      4@              I@      *@      �?      @              �?      �?      @      �?                      @     �H@       @      9@       @      2@       @      2@      @      1@      �?       @      �?      @              @      �?       @              �?      �?              �?      �?              "@              �?      @      �?      @              �?               @      @              8@                      @     �P@      @      1@             �H@      @      �?      �?      �?                      �?      H@       @      @       @      @                       @     �F@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJt�mUhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM=huh*h-K ��h/��R�(KM=��h|�B@O         ^                    �?�Qc�!�?�           @�@                                    @���!pc�?�            @n@                                   �?�-�[�?R            ``@                                  �?t�U����?,            �P@               
                    �?@4և���?             <@              	                 hލC@�t����?             1@                                `v7<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        
             ,@        ������������������������       �                     &@                                   �?8�Z$���?            �C@       ������������������������       �                     5@                                ���`@�q�q�?             2@       ������������������������       �                     "@                                    @�q�q�?             "@                               Ъ�c@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        &             P@               W                 ��Y7@�f��`��?H            �[@              P                    �?ƈ�VM�?9            @V@              ;                    ;@��S���?1            �R@              (                    1@8�A�0��?             F@                                ��,@���Q��?             4@        ������������������������       �                     @                                �L�@և���X�?             ,@        ������������������������       �                      @               #                    �?      �?             (@               "                    �?���Q��?             @               !                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        $       '                    @և���X�?             @       %       &                 P��%@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        )       2                 P�@      �?             8@        *       +                    �?����X�?             @        ������������������������       �                     �?        ,       -                 pf�@r�q��?             @        ������������������������       �                      @        .       1                 �&B@      �?             @       /       0                   �7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        3       4                  �#@�IєX�?
             1@        ������������������������       �                     &@        5       :                    �?r�q��?             @       6       9                    �?�q�q�?             @       7       8                    4@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        <       O                    B@¦	^_�?             ?@       =       H                    �?�+$�jP�?             ;@       >       ?                    �?�KM�]�?             3@        ������������������������       �                     @        @       A                 ���@r�q��?
             (@        ������������������������       �                     �?        B       G                    �?�C��2(�?	             &@       C       D                 ���@      �?              @        ������������������������       �                      @        E       F                 �&B@r�q��?             @       ������������������������       �      �?             @        ������������������������       �                      @        ������������������������       �                     @        I       L                 ��1@      �?              @       J       K                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        M       N                    3@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        Q       R                 ���&@؇���X�?             ,@        ������������������������       �                     �?        S       V                 ���.@$�q-�?             *@        T       U                   �<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        X       Y                    @���7�?             6@        ������������������������       �                     $@        Z       ]                    @�8��8��?             (@        [       \                 ��T?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        _       �                    �?z�G�z�?%           `}@        `       {                  I>@      �?)             P@       a       z                    �?ZՏ�m|�?            �H@       b       w                    �?��s����?             E@       c       l                    ;@8�Z$���?            �C@        d       e                 �{@      �?             @        ������������������������       �                     �?        f       g                 hfF&@���Q��?             @        ������������������������       �                      @        h       i                 ���0@�q�q�?             @        ������������������������       �                     �?        j       k                   �2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        m       v                 ���,@�C��2(�?            �@@       n       o                     @��2(&�?             6@        ������������������������       �                     �?        p       q                 ���@�����?             5@        ������������������������       �                      @        r       u                   @@8�Z$���?	             *@       s       t                    =@"pc�
�?             &@       ������������������������       ��<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     &@        x       y                @�µ2@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        |       �                   �;@��S���?             .@        }       �                   �7@z�G�z�?             @        ~                           �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?���Q��?             $@        �       �                    �?���Q��?             @       �       �                    >@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?z�G�z�?             @        ������������������������       �                     �?        �       �                   @K@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�@����?�            `y@        �       �                     @��� ��?             ?@        ������������������������       �                     @        �       �                   `3@؇���X�?             <@       �       �                    �?�C��2(�?             6@       �       �                  s�@�����?             5@        ������������������������       �                      @        �       �                    >@8�Z$���?             *@       �       �                   �<@z�G�z�?	             $@       �       �                 ��(@�����H�?             "@       ������������������������       �؇���X�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                     �?�.��7F�?�            pw@        �       �                   �J@t�C�#��?.            �S@       �       �                   �G@�G�z��?&             N@       �       �                     @���Q �?!            �H@       �       �                    �?r�qG�?              H@       �       �                   �E@v�X��?             F@       �       �                   �D@4�B��?            �B@       �       �                 `fF:@�������?             A@        ������������������������       �                     &@        �       �                   @B@�û��|�?             7@       �       �                    �?�q�q�?             2@       �       �                   �>@ҳ�wY;�?             1@        �       �                 `fF<@����X�?             @        ������������������������       ��q�q�?             @        ������������������������       �                     @        �       �                   �<@ףp=
�?	             $@       �       �                 ��yC@r�q��?             @        �       �                   �A@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �B@���Q��?             @        ������������������������       �                      @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �F@؇���X�?             @       �       �                    �?z�G�z�?             @       �       �                 `f?@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        �       �                   �R@�KM�]�?             3@       ������������������������       �                     1@        ������������������������       �                      @        �       �                    @���G��?�            �r@        �       �                    �?     ��?
             0@       �       �                   �C@����X�?             ,@       �       �                     @r�q��?             (@       ������������������������       �                     @        �       �                    @���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       <                  @E@$s��O�?�            �q@       �       9                  �D@L�S5]�?�             n@       �       8                   �?��E�B��?�            `m@       �       1                0��D@�{�9�?�            `j@       �       0                   �?pLBQh��?�             i@       �       �                 @33@0sS]�?~            �h@        �       �                   �:@X�<ݚ�?             "@        �       �                    6@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 �?�@p�/E�f�?y            �g@        �       �                   �4@@4և���?0             U@        ������������������������       �        	             3@        �       �                 pb@���Ls�?'            @P@       �       �                 �?$@�p ��?            �D@       �       �                    �?l��\��?             A@       �       �                 ���@�C��2(�?            �@@        ������������������������       �                     $@        �       �                 ���@�LQ�1	�?             7@        ������������������������       �                      @        �       �                 ���@���N8�?             5@       ������������������������       �                     ,@        �       �                   �=@؇���X�?             @        �       �                    ;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �5@և���X�?             @        ������������������������       �                      @        �       �                   �9@z�G�z�?             @        ������������������������       �                     @        �       �                   �;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     8@        �                       @3�@T�6|���?I             Z@        �                          �?      �?              @       �                         �A@����X�?             @       �                         �?@r�q��?             @                                  :@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?              )                   �?      �?C             X@                               �<@���H��?<             U@                                 @6uH���?,             O@        	                         &@$�q-�?             :@        
                        �5@؇���X�?             @                               �1@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     @                                �;@�}�+r��?             3@       ������������������������       �                     0@                                �*@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                              @�!@�8��8��?             B@                             ��) @�LQ�1	�?             7@                               �3@@4և���?
             ,@        ������������������������       �                     �?        ������������������������       �        	             *@                                �7@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        	             *@              $                  @@@�GN�z�?             6@              #                   $@���Q��?             $@              "                  �>@z�G�z�?             @              !                �̌!@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        %      (                  @A@�8��8��?
             (@        &      '                    @z�G�z�?             @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     @        *      +                м�6@r�q��?             (@       ������������������������       �                     @        ,      /                  �@@�q�q�?             @       -      .                  �<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        2      3                    @      �?             $@        ������������������������       �                      @        4      5                   ;@      �?              @        ������������������������       �                      @        6      7                   >@      �?             @       ������������������������       �      �?             @        ������������������������       �                      @        ������������������������       �                     8@        :      ;                   �?�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                    �C@        �t�bh�h*h-K ��h/��R�(KM=KK��h]�B�       �{@     �p@     �P@      f@       @     �^@       @     �M@       @      :@       @      .@       @      �?              �?       @                      ,@              &@      @     �@@              5@      @      (@              "@      @      @      @      �?      @                      �?               @              P@      M@     �J@     �B@      J@     �A@      D@      :@      2@       @      (@              @       @      @       @              @      @       @      @       @      �?       @                      �?               @      @      @       @      @       @                      @       @              2@      @       @      @      �?              �?      @               @      �?      @      �?      �?              �?      �?                       @      0@      �?      &@              @      �?       @      �?      �?      �?              �?      �?              �?              @              "@      6@      @      6@       @      1@              @       @      $@      �?              �?      $@      �?      @               @      �?      @      �?      @               @              @      @      @      �?      @              @      �?               @      �?       @                      �?      @               @      (@      �?              �?      (@      �?       @      �?                       @              $@      5@      �?      $@              &@      �?      �?      �?      �?                      �?      $@             �w@     �W@      H@      0@     �D@       @      A@       @     �@@      @      @      @      �?               @      @               @       @      �?      �?              �?      �?      �?                      �?      >@      @      3@      @              �?      3@       @       @              &@       @      "@       @      @       @       @               @              &@              �?       @               @      �?              @              @       @      �?      @      �?      �?      �?                      �?              @      @      @       @      @       @      �?       @                      �?               @      @      �?      �?              @      �?      @                      �?     �t@     �S@      ;@      @      @              8@      @      4@       @      3@       @       @              &@       @       @       @       @      �?      @      �?       @                      �?      @              �?              @       @      @                       @     �r@     �R@      I@      =@     �@@      ;@      @@      1@      ?@      1@      ?@      *@      9@      (@      9@      "@      &@              ,@      "@      (@      @      &@      @       @      @       @      �?              @      "@      �?      @      �?       @      �?       @                      �?      @              @              �?               @      @               @       @      �?       @                      �?              @      @      �?      @      �?       @      �?      �?      �?      �?               @               @                      @      �?              �?      $@              $@      �?              1@       @      1@                       @     `o@     �F@      @      &@      @      $@       @      $@              @       @      @       @                      @       @              �?      �?              �?      �?             �n@      A@     �i@      A@     �i@      >@     �f@      >@      f@      9@     �e@      9@      @      @      �?      @      �?                      @      @             �d@      5@     �S@      @      3@             �M@      @     �A@      @      ?@      @      >@      @      $@              4@      @               @      4@      �?      ,@              @      �?      �?      �?      �?                      �?      @              �?              @      @               @      @      �?      @              �?      �?              �?      �?              8@             @V@      .@      @      @      @       @      @      �?      �?      �?      �?                      �?      @                      �?              �?      U@      (@     �R@      $@     �L@      @      8@       @      @      �?      @      �?      �?               @      �?      @              2@      �?      0@               @      �?              �?       @             �@@      @      4@      @      *@      �?              �?      *@              @       @      @                       @      *@              1@      @      @      @      �?      @      �?       @      �?                       @               @      @              &@      �?      @      �?      �?      �?      @              @              $@       @      @              @       @      �?       @      �?                       @      @              @              @      @       @              @      @               @      @      @      @      �?               @      8@               @      @              @       @             �C@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJc��hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM/huh*h-K ��h/��R�(KM/��h|�B�K                             �?�uY0�l�?�           @�@                                   @�����H�?	             "@       ������������������������       �                      @        ������������������������       �                     �?               X                     �?6�t��?�           ��@               5                   �D@���a���?j            �d@                                `fK@θ	j*�?C             Z@               	                    �?�q�q�?             ;@        ������������������������       �                     @        
                           B@      �?             8@                                  �?����X�?             5@                                  �?     ��?             0@        ������������������������       �                     �?                                   @@������?             .@                                 �<@d}h���?             ,@                               ��yC@�θ�?
             *@                               `fF:@�q�q�?             "@        ������������������������       �                     @                                `f�<@      �?             @        ������������������������       �                      @                                  �A@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?                                `fFJ@z�G�z�?             @        ������������������������       �                     @                                   7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        !       $                    �?6��f�?0            @S@       "       #                     @p���?             I@        ������������������������       �                     �?        ������������������������       �                    �H@        %       0                    >@X�<ݚ�?             ;@       &       -                    �?�E��ӭ�?             2@       '       (                   �1@���|���?             &@        ������������������������       �                     �?        )       ,                    �?�z�G��?             $@       *       +                 ���S@      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        .       /                    '@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        1       4                    �?�<ݚ�?             "@        2       3                 pU�t@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        6       W                 ��^@�^�����?'             O@       7       >                    �?>4և���?#             L@        8       9                   �H@�KM�]�?             3@        ������������������������       �                     $@        :       =                 83F@�<ݚ�?             "@        ;       <                 ���;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ?       V                   �R@�MI8d�?            �B@       @       M                    �?(N:!���?            �A@        A       F                    �?���!pc�?             &@        B       E                   �L@      �?             @       C       D                   �I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        G       H                   @H@����X�?             @        ������������������������       �                     �?        I       L                    �?r�q��?             @       J       K                 @�pX@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        N       O                    �? �q�q�?             8@        ������������������������       �                      @        P       U                 `f�;@���7�?             6@        Q       T                    J@�C��2(�?             &@        R       S                   �G@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             &@        ������������������������       �                      @        ������������������������       �                     @        Y       �                 `f�$@f��kG|�?R           Ȁ@        Z       �                   @@@LH=$��?�            Pp@       [       x                    �?�!�z�0�?�            �j@        \       m                  ��@��S���?             �F@       ]       ^                 03�@�q�q�?             8@        ������������������������       �                     �?        _       f                 ���@�㙢�c�?             7@       `       a                    �?$�q-�?	             *@        ������������������������       �                     @        b       e                 ���@�����H�?             "@        c       d                    9@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        g       h                   �9@�z�G��?             $@        ������������������������       �                      @        i       j                    ;@      �?              @        ������������������������       �                      @        k       l                 �&B@r�q��?             @       ������������������������       ��q�q�?             @        ������������������������       �                     @        n       q                    �?���N8�?             5@        o       p                   �5@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        r       w                   �>@���y4F�?             3@       s       v                   �2@      �?             0@        t       u                     @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             ,@        ������������������������       �                     @        y       z                     @$�Q�\�?i             e@        ������������������������       �                     @        {       �                   �?@�<p���?g            �d@       |       �                   �;@X��P�T�?c            �c@        }       �                    �?���!���?0            �S@        ~                        ���@�q�q�?             @        ������������������������       �                     �?        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�KM�]�?-             S@       �       �                 �1@�����H�?+             R@        �       �                    7@tk~X��?             B@       �       �                 �?$@ �q�q�?             8@       ������������������������       �        	             6@        �       �                   �5@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?      �?             (@        ������������������������       �                      @        �       �                 �&b@���Q��?             $@        �       �                 @33@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    9@r�q��?             @        ������������������������       �                     @        �       �                   �:@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �0@������?             B@        ������������������������       �      �?              @        ������������������������       �                     A@        ������������������������       �                     @        �       �                 ���"@ �\���?3            �S@       �       �                 ��@xL��N�?0            �R@        �       �                   @<@�#-���?            �A@       �       �                 ���@ �Cc}�?             <@        ������������������������       �                     @        �       �                 �Y�@؇���X�?             5@        ������������������������       ����Q��?             @        �       �                    �?      �?
             0@       �       �                  s�@@4և���?             ,@        ������������������������       �                     @        �       �                    �?�C��2(�?             &@       ������������������������       ������H�?             "@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                    �C@        �       �                   �<@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 P�@r�q��?             @        ������������������������       �                      @        �       �                 @3�@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        �       �                 `f#@`Ql�R�?            �G@       ������������������������       �                     G@        ������������������������       �                     �?        �       $                   @�)
;&��?�            @q@       �       �                    @Z�K�D��?�            `m@        ������������������������       �                     @        �       �                    �?�LQ�1	�?�            �l@       �       �                    �?��w��?Q            ``@        �       �                    �?�חF�P�?             ?@        �       �                 ��	-@      �?             @        ������������������������       �                     �?        �       �                  S�2@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 @3�2@�����H�?             ;@       �       �                     @�}�+r��?             3@       �       �                    �?$�q-�?             *@        ������������������������       �                     �?        �       �                 `f�)@�8��8��?             (@        ������������������������       �                     @        �       �                    :@�����H�?             "@        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                 039@      �?              @        �       �                     @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                 0��D@0w-!��?8             Y@       �       �                   �4@��r
'��?4            @W@       �       �                 ��q1@�ݜ�?+            �S@       �       �                     @����1�?)            @R@       �       �                    �?Xny��?"            �N@        �       �                 `��,@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    &@ �Cc}�?             L@        �       �                   �H@d}h���?	             ,@       �       �                   �6@�C��2(�?             &@        �       �                   �1@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        �       �                   �P@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �*@@4և���?             E@       �       �                 `f�)@l��\��?             A@        ������������������������       �                     @        �       �                   �;@�����H�?             ;@        ������������������������       �                     $@        �       �                    =@@�0�!��?	             1@        ������������������������       �                     �?        �       �                    @@      �?             0@        ������������������������       �                     @        �       �                   @B@r�q��?             (@        ������������������������       �      �?             @        �       �                   @D@      �?              @        ������������������������       �                      @        �       �                   �G@r�q��?             @       ������������������������       �z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     (@        �       �                   �2@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        	             .@        �       �                 ��?P@և���X�?             @       �       �                    >@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                  s�+@F߼�q�?=            �X@        ������������������������       �                     @        �                          �?֭��F?�?;            �W@       �       
                  �;@f�Sc��?            �H@               	                  �H@      �?	             0@                                 @z�G�z�?             .@                                �3@      �?             @        ������������������������       �                      @        ������������������������       �                      @                              @3�/@�C��2(�?             &@                                 �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?                                  @"pc�
�?            �@@        ������������������������       �                     *@                              ��Y7@�z�G��?             4@                                �?      �?	             0@        ������������������������       �                     @                              ���.@z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @                                 �?�����H�?            �F@                                 @      �?             @@                              0C�:@�����H�?
             2@                               �@@"pc�
�?             &@                                �?���Q��?             @        ������������������������       �                     �?                                �>@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        
             ,@               #                `f62@�θ�?	             *@        !      "                �=/@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        %      .                  �>@������?            �D@       &      '                   �?�(\����?             D@        ������������������������       �                     &@        (      )                ��T?@XB���?             =@        ������������������������       �                     ,@        *      -                   @��S�ۿ?	             .@        +      ,                   @      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     �?        �t�bh�h*h-K ��h/��R�(KM/KK��h]�B�       �}@     �m@      �?       @               @      �?             �}@     �l@     �P@     �X@      A@     �Q@      2@      "@              @      2@      @      .@      @      &@      @              �?      &@      @      &@      @      $@      @      @      @      @              @      @               @      @      �?      @                      �?      @              �?                      �?      @      �?      @              �?      �?      �?                      �?      @              0@     �N@      �?     �H@      �?                     �H@      .@      (@      *@      @      @      @              �?      @      @      @      @              @      @               @              @      �?              �?      @               @      @       @      @       @                      @              @     �@@      =@     �@@      7@       @      1@              $@       @      @       @      �?              �?       @                      @      ?@      @      ?@      @       @      @      @      �?      �?      �?      �?                      �?       @              @       @              �?      @      �?       @      �?              �?       @              @              7@      �?       @              5@      �?      $@      �?      @      �?      @                      �?      @              &@                       @              @     py@     @`@     @k@     �E@     �e@      E@      5@      8@      @      3@      �?              @      3@      �?      (@              @      �?       @      �?       @               @      �?                      @      @      @       @              �?      @               @      �?      @      �?       @              @      0@      @      �?      �?              �?      �?              .@      @      .@      �?      �?      �?      �?                      �?      ,@                      @     �b@      2@      @             @b@      2@      b@      *@     �Q@      "@       @      �?      �?              �?      �?              �?      �?              Q@       @      P@       @      =@      @      7@      �?      6@              �?      �?              �?      �?              @      @       @              @      @      @      �?              �?      @              �?      @              @      �?       @      �?                       @     �A@      �?      �?      �?      A@              @             �R@      @     �Q@      @      @@      @      9@      @      @              2@      @      @       @      .@      �?      *@      �?      @              $@      �?       @      �?       @               @              @             �C@              @      �?      @                      �?      �?      @               @      �?      @      �?       @              �?      G@      �?      G@                      �?     �g@     �U@     �b@     @U@              @     �b@      T@      W@     �C@      @      :@       @       @              �?       @      �?       @                      �?      @      8@      �?      2@      �?      (@              �?      �?      &@              @      �?       @      �?       @              @              @       @      @       @      �?              �?       @                      @     �U@      *@     �T@      $@      Q@      $@     �P@      @      K@      @      @      �?              �?      @              I@      @      &@      @      $@      �?      �?      �?      �?                      �?      "@              �?       @               @      �?             �C@      @      ?@      @      @              8@      @      $@              ,@      @              �?      ,@       @      @              $@       @      @      �?      @      �?       @              @      �?      @      �?      �?               @              (@               @      @       @                      @      .@              @      @       @      @       @                      @       @              M@     �D@              @      M@      B@      2@      ?@      (@      @      (@      @       @       @               @       @              $@      �?       @      �?       @                      �?       @                      �?      @      ;@              *@      @      ,@       @      ,@              @       @       @       @                       @      @              D@      @      >@       @      0@       @      "@       @      @       @      �?               @       @       @                       @      @              @              ,@              $@      @      @      @      @                      @      @             �C@       @     �C@      �?      &@              <@      �?      ,@              ,@      �?      @      �?      @                      �?      &@                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJg�$hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM#huh*h-K ��h/��R�(KM#��h|�B�H         b                    �?(����7�?�           @�@               a                    @0,Tg��?�            �o@              `                    @���?�            �n@              %                     @�mEx���?�             n@                                   �?0Ƭ!sĮ?Y             `@                                  �?Pa�	�?0            �P@                                   �?h�����?             <@                                  �?P���Q�?             4@       	       
                   �G@�X�<ݺ?             2@       ������������������������       �        	             ,@                                ,w�U@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @                                   �?P�Lt�<�?             C@        ������������������������       �                     6@                                   �?      �?             0@       ������������������������       �        
             (@                                  �8@      �?             @        ������������������������       �                      @                                  �>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               $                   �;@�i�y�?)            �O@                                  �?�>����?             ;@        ������������������������       �                     "@               #                    �?�����H�?             2@                                    �?�q�q�?             @                                 �6@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        !       "                    7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                     B@        &       ;                    �?������?>             \@        '       :                 ��.@�t����?            �I@       (       9                    �?��]�T��?            �D@       )       8                 P��+@�E��ӭ�?             B@       *       /                 ���@     ��?             @@        +       ,                   �5@      �?              @        ������������������������       �                      @        -       .                 0��@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        0       7                    �?�8��8��?             8@       1       4                   �5@���}<S�?             7@        2       3                    2@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        5       6                 pF @�}�+r��?
             3@       ������������������������       �        	             2@        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@        <       [                    �?Nd^����?#            �N@       =       L                   �;@�û��|�?             G@       >       I                    �?և���X�?             5@       ?       @                   �4@      �?             0@        ������������������������       �                     @        A       H                    �?�θ�?             *@       B       G                 03�!@���!pc�?             &@       C       D                   �7@�����H�?             "@        ������������������������       �                     @        E       F                 �&B@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        J       K                   �8@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        M       X                    �?�+e�X�?             9@       N       O                 03�!@������?             .@        ������������������������       �                     @        P       W                 ��1@X�<ݚ�?             "@       Q       V                    �?�q�q�?             @       R       U                   &@      �?             @       S       T                    I@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        Y       Z                   �>@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        \       ]                 �̼6@��S���?             .@        ������������������������       �                     @        ^       _                    @���!pc�?             &@       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        c       r                    *@�܆!�t�?"           �|@        d       i                    �?�q�q�?             8@        e       f                    @؇���X�?             @        ������������������������       �                     @        g       h                 �y.@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        j       q                    $@j���� �?             1@       k       l                    @      �?             0@        ������������������������       �                     "@        m       n                 ��A>@؇���X�?             @        ������������������������       �                     @        o       p                 ���A@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        s       �                    �?��UTF@�?           @{@        t       �                 xCQ@�n_Y�K�?,            �S@       u       �                    ;@�<ݚ�?"             K@        v       w                   �1@�z�G��?             $@        ������������������������       �                     �?        x                           �?�<ݚ�?             "@       y       ~                    �?      �?              @       z       {                 ���@z�G�z�?             @        ������������������������       �                     @        |       }                    8@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �J@�Ra����?             F@       �       �                    �?$�q-�?            �C@       �       �                    �?l��\��?             A@       �       �                   @@@ףp=
�?             >@       �       �                   �<@�S����?             3@       �       �                     �?�IєX�?             1@        �       �                 03SA@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        
             ,@        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �                     @        ������������������������       �                     @        �       �                 ��L@@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?      �?
             8@       �       �                 @�?t@�q�q�?             2@       �       �                   �8@      �?             (@        ������������������������       �                     @        �       �                   @B@�q�q�?             "@        ������������������������       �                     @        �       �                  �}S@      �?             @        ������������������������       �                      @        �       �                   �G@      �?             @        ������������������������       �                      @        �       �                   �H@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 `ff:@@�qmNh�?�            `v@       �       �                   @@@��� =�?�             q@       �       �                 ��@�^'�ë�?�            @h@        �       �                   �;@ �#�Ѵ�?            �E@        �       �                    @؇���X�?             ,@        ������������������������       �                     �?        �       �                    �?$�q-�?
             *@        ������������������������       �                     @        �       �                 ��@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     =@        �       �                   �>@*~k���?e            �b@       �       �                    �?�1�hP	�?^            �a@       �       �                   �4@�u����?Z             a@        �       �                     @z�G�z�?            �A@        �       �                    &@�q�q�?             "@        �       �                   �1@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   �0@8�Z$���?             :@        �       �                 �̌!@����X�?             @       �       �                 pf�@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     @        �       �                    �?�KM�]�?             3@       �       �                 ��Y @�X�<ݺ?             2@       �       �                 �?�@ףp=
�?             $@       ������������������������       �                     @        �       �                   �3@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                 �?$@�:�]��?C            �Y@        ������������������������       �                      @        �       �                    �? "��u�?A             Y@        �       �                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�}�+r��?>            �W@       �       �                   �:@ ��Ou��?2            �S@        ������������������������       �                    �A@        �       �                     @X�EQ]N�?            �E@        �       �                   �3@؇���X�?             @       �       �                   �<@z�G�z�?             @        �       �                   �;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                 ��) @�����H�?             B@       �       �                   �;@ ��WV�?             :@        ������������������������       �                     �?        ������������������������       �                     9@        �       �                   �;@�z�G��?             $@        ������������������������       �                     �?        �       �                 pf� @�<ݚ�?             "@        ������������������������       �                     �?        �       �                 ��)"@      �?              @        ������������������������       �                      @        �       �                   �<@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     1@        ������������������������       �                     @        �       �                     @      �?              @        ������������������������       �                     �?        �       �                    �?����X�?             @       �       �                   �?@���Q��?             @        ������������������������       �                     �?        �       �                   �@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�(�Tw�?2            �S@       �       �                 @3�@@	tbA@�?,            @Q@        �       �                   �B@�nkK�?             7@        ������������������������       �                     $@        �       �                    �?$�q-�?             *@        ������������������������       �                     �?        �       �                      @�8��8��?
             (@        ������������������������       �                     @        �       �                 �?�@�����H�?             "@       ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     G@        ������������������������       �                     "@        �                         �>@p����?1            �U@        �                          �?�G��l��?             5@       �                          L@      �?             4@       �                         @G@�q�q�?             .@       �                           �?X�<ݚ�?             "@                                @B@      �?              @                             `fF<@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        	                         �?��ɉ�?%            @P@       
                         �?z�G�z�?             D@        ������������������������       �                     �?                                 D@x�����?            �C@                                �?r֛w���?             ?@                                �?����X�?             <@                               �?@�z�G��?             4@                                 @�<ݚ�?
             2@       ������������������������       �                     (@                                 ;@�q�q�?             @        ������������������������       �                      @        ������������������������       �      �?             @        ������������������������       �                      @                              03U@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @              "                    �?`2U0*��?             9@                                �?�8��8��?             (@        ������������������������       �                     @              !                    @�����H�?             "@                               x�N@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     *@        �t�b��     h�h*h-K ��h/��R�(KM#KK��h]�B0       �{@      q@     �P@     @g@      N@     @g@     �K@     @g@      @     @_@       @      P@      �?      ;@      �?      3@      �?      1@              ,@      �?      @      �?                      @               @               @      �?     �B@              6@      �?      .@              (@      �?      @               @      �?      �?      �?                      �?       @     �N@       @      9@              "@       @      0@       @      @      �?      @              �?      �?       @      �?      �?              �?      �?                      (@              B@     �I@     �N@      .@      B@      .@      :@      $@      :@      @      :@      @      @               @      @       @               @      @               @      6@       @      5@      �?      @              @      �?              �?      2@              2@      �?                      �?      @              @                      $@      B@      9@      <@      2@      "@      (@      @      $@      @              @      $@      @       @      �?       @              @      �?      @      �?                      @       @                       @      @       @               @      @              3@      @      &@      @      @              @      @       @      @       @       @       @      �?       @                      �?              �?               @      @               @       @       @                       @       @      @              @       @      @       @                      @      @              @             `w@     �U@       @      0@      �?      @              @      �?      @              @      �?              @      $@      @      $@              "@      @      �?      @               @      �?              �?       @              �?             �v@     �Q@      H@      >@      E@      (@      @      @      �?               @      @      �?      @      �?      @              @      �?      �?      �?                      �?              @      �?             �C@      @      B@      @      ?@      @      ;@      @      0@      @      0@      �?       @      �?              �?       @              ,@                       @      &@              @              @              @       @      @                       @      @      2@      @      (@      @      @      @              @      @              @      @      @               @      @      �?       @              �?      �?              �?      �?                      @              @     �s@      D@     `o@      5@     �e@      4@     �D@       @      (@       @              �?      (@      �?      @               @      �?              �?       @              =@             �`@      2@      `@      .@     �^@      .@      <@      @      @      @      �?      @      �?                      @      @              6@      @      @       @       @       @      �?              �?       @      @              1@       @      1@      �?      "@      �?      @               @      �?      �?      �?      �?               @                      �?     �W@       @               @     �W@      @      @      �?      @                      �?     �V@      @     @R@      @     �A@              C@      @      @      �?      @      �?      �?      �?      �?                      �?      @               @              @@      @      9@      �?              �?      9@              @      @              �?      @       @              �?      @      �?       @              @      �?      @                      �?      1@              @              @      @              �?      @       @      @       @              �?      @      �?              �?      @               @             @S@      �?      Q@      �?      6@      �?      $@              (@      �?      �?              &@      �?      @               @      �?      @              �?      �?      G@              "@             �P@      3@      &@      $@      $@      $@      @      $@      @      @      @      @      �?      @      �?                      @      @              �?                      @      @              �?              L@      "@      @@       @      �?              ?@       @      7@       @      4@       @      ,@      @      ,@      @      (@               @      @               @       @       @               @      @       @      @                       @      @               @              8@      �?      &@      �?      @               @      �?      @      �?              �?      @               @              *@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�>D5hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM'huh*h-K ��h/��R�(KM'��h|�B�I                             @Dl���v�?�           @�@                                   @��<b���?             G@                               P��%@г�wY;�?             A@                                �(\�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @@               	                 ��T?@      �?             (@        ������������������������       �                     @        
                        ���A@      �?             @        ������������������������       �                     @        ������������������������       �                     @               f                    �?D��J<��?�           Є@               U                    �?��eN_:�?�             j@              "                     @B�0�~d�?w             f@                               03�a@ 5x ��?E            �Z@                                  �?�q�q�??             X@                                �v7@0�z��?�?.             O@                                   �?P���Q�?             4@        ������������������������       �                     @                                  �;@�IєX�?             1@                                   8@      �?             @        ������������������������       �                     �?                                  �/@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        
             *@        ������������������������       �                     E@        ������������������������       �                     A@                                   �?"pc�
�?             &@       ������������������������       �                      @                !                   �A@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        #       B                    �?������?2            @Q@       $       =                    �?�û��|�?!             G@       %       <                    �?#z�i��?            �D@       &       '                    �?p�ݯ��?             C@        ������������������������       �                     @        (       )                   �5@j���� �?             A@        ������������������������       �                     @        *       1                 �̌@8^s]e�?             =@       +       0                   @B@�����H�?             2@       ,       /                 ���@�IєX�?             1@        -       .                    9@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        
             .@        ������������������������       �                     �?        2       ;                   @G@���|���?             &@       3       :                 @3S%@�<ݚ�?             "@       4       5                    �?      �?              @        ������������������������       �                     �?        6       9                 @3�@؇���X�?             @        7       8                 �?�@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        >       ?                  S�2@z�G�z�?             @        ������������������������       �                     @        @       A                 �A7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        C       T                   �B@�û��|�?             7@       D       Q                    �?�\��N��?             3@       E       L                    ;@��S���?             .@        F       K                   �8@r�q��?             @       G       H                    �?�q�q�?             @        ������������������������       �                     �?        I       J                    6@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        M       N                   �=@�<ݚ�?             "@       ������������������������       �                     @        O       P                   �@@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        R       S                   @@@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        V       W                   �0@�eP*L��?            �@@        ������������������������       �                     @        X       e                    @
j*D>�?             :@       Y       d                    =@      �?             8@       Z       c                   �b@�\��N��?
             3@       [       \                    �?X�Cc�?             ,@        ������������������������       �                      @        ]       b                 м6@      �?             (@        ^       _                   �1@      �?             @        ������������������������       �                      @        `       a                    5@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        g       &                   @���2���?!           �|@       h       �                   �<@>.��Y��?           `|@       i       x                   �1@*
;&���?�            @q@        j       w                    @     ��?             @@       k       l                    $@      �?             6@        ������������������������       �                     @        m       v                    �?D�n�3�?             3@       n       u                    �?     ��?             0@       o       r                 pf� @X�Cc�?             ,@        p       q                 pf�@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        s       t                    �?�����H�?	             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     $@        y       �                 �?$@�&�4rd�?�            �n@        z       {                 ���@"pc�
�?.             V@        ������������������������       �                     ,@        |       }                 ��@���@��?&            �R@        ������������������������       �                     @        ~       �                   �9@O�o9%�?%            �Q@               �                 �Y�@R�}e�.�?             :@        �       �                 ���@      �?             (@        ������������������������       �                     @        �       �                    5@؇���X�?             @        ������������������������       �                      @        �       �                    �?z�G�z�?             @       �       �                 ���@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ��@@4և���?             ,@       ������������������������       �                     "@        �       �                    �?z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�r����?            �F@       �       �                   @<@��2(&�?             F@       �       �                    ;@؇���X�?             E@        ������������������������       �                     �?        �       �                    �?�p ��?            �D@       �       �                 ���@HP�s��?
             9@        ������������������������       �                     &@        ������������������������       �؇���X�?             ,@        �       �                 ��@      �?	             0@       �       �                    �?z�G�z�?             .@       �       �                  s�@���!pc�?             &@        ������������������������       �                      @        ������������������������       ��q�q�?             "@        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                     �?4��?�?f            �c@        �       �                   �8@r֛w���?             ?@        ������������������������       �                     $@        �       �                    �?�ՙ/�?             5@        �       �                   �;@���!pc�?             &@        �       �                 hD�b@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?      �?             $@       �       �                 ��9B@X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?@�E~��?P            @_@        �       �                 033.@���!pc�?             &@       ������������������������       �                     @        �       �                   �6@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?���U�?J            �\@        �       �                   `3@      �?              @       ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �*@�|1)�?E            �Z@       �       �                     @`2U0*��?3            �R@        �       �                   �;@P���Q�?             4@       ������������������������       �        	             2@        �       �                   �'@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �3@h㱪��?(            �K@        �       �                   �2@؇���X�?             @        ������������������������       �                     @        �       �                 `�8"@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        �       �                 ��) @@��8��?#             H@       ������������������������       �                    �C@        �       �                 pf� @�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     ?@        �       %                ��M\@�μ���?v            @f@       �                        ��$:@��q���?r            `e@       �       �                   �=@>4և�z�?K             \@        �       �                    �?�q�q�?             "@        ������������������������       �                     @        �       �                    $@      �?             @       �       �                 �̌!@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   �F@���z�k�?F            �Y@       �       �                    �?�?�'�@�?0             S@       �       �                     @8�Z$���?+            @P@        �       �                    1@�θ�?             *@       �       �                     �?      �?              @        ������������������������       �                     �?        �       �                    @@և���X�?             @        ������������������������       �                      @        ������������������������       ����Q��?             @        ������������������������       �                     @        �       �                 �?�@���c���?              J@        �       �                   @@@ 7���B�?             ;@        �       �                 �&B@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             5@        �       �                    �?�+e�X�?             9@       �       �                 @3�@����X�?             5@        �       �                   �D@      �?              @       �       �                   �?@���Q��?             @        ������������������������       �                     �?        �       �                   �A@      �?             @        ������������������������       �                      @        ������������������������       �      �?              @        ������������������������       �                     @        �       �                 ��i @$�q-�?
             *@       �       �                   �@@      �?              @        �       �                    ?@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     &@        �       �                    �? 7���B�?             ;@        ������������������������       �                      @        �       �                 `f'@`2U0*��?             9@       �       �                   �#@$�q-�?             *@       ������������������������       �        	             &@        �       �                   �P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             (@                              03k:@L
�q��?'            �M@        ������������������������       �                     @                                �?@Dc}h��?&             L@        ������������������������       �                      @                                 �?r�qG�?"             H@                                 �?և���X�?	             ,@                               �H@�q�q�?             (@                               �G@�z�G��?             $@       	      
                   A@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @                                 �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?              $                    @�������?             A@             #                   �?r٣����?            �@@             "                03�U@����X�?             <@                                @@������?             ;@                               @=@      �?             0@                             `f�;@����X�?
             ,@                               �J@�	j*D�?	             *@                                @G@z�G�z�?             @        ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @              !                  �C@�C��2(�?	             &@                                  �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �t�bh�h*h-K ��h/��R�(KM'KK��h]�Bp        {@     `q@      $@      B@      �?     �@@      �?      �?              �?      �?                      @@      "@      @      @              @      @              @      @             �z@     @n@     �J@     �c@     �A@     �a@      @      Z@      �?     �W@      �?     �N@      �?      3@              @      �?      0@      �?      @              �?      �?       @               @      �?                      *@              E@              A@       @      "@               @       @      �?       @                      �?      @@     �B@      2@      <@      ,@      ;@      ,@      8@              @      ,@      4@      @              "@      4@       @      0@      �?      0@      �?      �?              �?      �?                      .@      �?              @      @      @       @      @      �?      �?              @      �?       @      �?       @                      �?      @                      �?               @              @      @      �?      @              �?      �?              �?      �?              ,@      "@      $@      "@      @       @      @      �?       @      �?      �?              �?      �?      �?                      �?      @               @      @              @       @      �?       @                      �?      @      �?      @                      �?      @              2@      .@      @              &@      .@      "@      .@      "@      $@      "@      @               @      "@      @      �?      @               @      �?      �?      �?                      �?       @                      @              @       @             0w@     �U@      w@     �U@     @m@      E@      5@      &@      &@      &@              @      &@       @      &@      @      "@      @      �?      @      �?                      @       @      �?       @                      �?       @                      @      $@             �j@      ?@      R@      0@      ,@              M@      0@              @      M@      *@      3@      @      @      @      @              �?      @               @      �?      @      �?      @              @      �?                      �?      *@      �?      "@              @      �?      @                      �?     �C@      @      C@      @      B@      @      �?             �A@      @      7@       @      &@              (@       @      (@      @      (@      @       @      @       @              @      @      @                      �?       @              �?             �a@      .@      7@       @      $@              *@       @       @      @      �?      @              @      �?              @              @      @      @      @              @      @                      �?     �]@      @       @      @      @              �?      @              @      �?             �[@      @      @      �?      @               @      �?       @                      �?     �Y@      @      R@      @      3@      �?      2@              �?      �?      �?                      �?     �J@       @      @      �?      @              @      �?       @      �?      �?             �G@      �?     �C@               @      �?              �?       @              ?@             �`@      F@     �`@     �B@     �W@      1@      @      @              @      @      @      �?      @      �?                      @       @              W@      &@     �P@      $@     �K@      $@      $@      @      @      @      �?              @      @       @               @      @      @             �F@      @      :@      �?      @      �?      @                      �?      5@              3@      @      .@      @      @      @      @       @              �?      @      �?       @              �?      �?              @      (@      �?      @      �?       @      �?       @                      �?      @              @              @              &@              :@      �?       @              8@      �?      (@      �?      &@              �?      �?              �?      �?              (@             �C@      4@              @     �C@      1@       @              ?@      1@      @       @      @      @      @      @      @       @               @      @                      @       @              �?      �?      �?                      �?      9@      "@      9@       @      4@       @      4@      @      $@      @      $@      @      "@      @      �?      @      �?       @               @       @              �?                       @      $@      �?       @      �?       @                      �?       @                      �?      @                      �?              @      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ���&hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM%huh*h-K ��h/��R�(KM%��h|�B@I         b                    �?T�����?�           @�@                                    @^������?�            �n@                                  �?P���Q�?P             ^@                                   �?����D��?A            @W@       ������������������������       �        %            �I@                                   �?���N8�?             E@       ������������������������       �                     =@                                   �?8�Z$���?             *@       	                           �?      �?              @       
                           �?���Q��?             @        ������������������������       �                      @                                  �9@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @                                   �?PN��T'�?             ;@        ������������������������       �                     &@                                ���`@      �?
             0@       ������������������������       �                     "@                                   �?և���X�?             @        ������������������������       �                     @        ������������������������       �                     @               E                    �?z�m�(�?D            @_@              2                    �?��:c���?'            �P@                                03�@      �?             @@        ������������������������       �                     @               +                    �?П[;U��?             =@                                  �?�t����?             1@        ������������������������       �                     @                                 ���@�n_Y�K�?
             *@        ������������������������       �                      @        !       $                   �5@���!pc�?	             &@        "       #                  s�@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        %       &                    9@�<ݚ�?             "@        ������������������������       �                      @        '       (                 ���@����X�?             @        ������������������������       �                      @        )       *                 �&B@���Q��?             @        ������������������������       ��q�q�?             @        ������������������������       �                      @        ,       -                 03�-@�q�q�?             (@        ������������������������       �                     @        .       1                   �<@      �?              @       /       0                    -@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        3       @                   �;@���Q��?            �A@       4       5                 ���@
;&����?             7@        ������������������������       �                     @        6       ?                   �9@b�2�tk�?             2@       7       >                 ��)+@d}h���?             ,@       8       =                    4@�8��8��?             (@        9       :                 x&�!@z�G�z�?             @        ������������������������       �                      @        ;       <                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        A       B                 `�X!@r�q��?             (@        ������������������������       �                     @        C       D                    >@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        F       ]                    �?����S��?             M@       G       H                    @�Gi����?            �B@        ������������������������       �                     @        I       Z                    @�q�q�?            �@@       J       U                    �?X�Cc�?             <@       K       L                   �6@�E��ӭ�?             2@        ������������������������       �                     @        M       T                    �?�q�q�?             (@       N       O                    �?���|���?             &@        ������������������������       �                     @        P       Q                    �?և���X�?             @        ������������������������       �                     �?        R       S                 @3S)@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        V       Y                   �>@      �?             $@       W       X                    �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        [       \                   �>@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ^       _                 ��T?@�����?	             5@       ������������������������       �                     *@        `       a                    @      �?              @        ������������������������       �                      @        ������������������������       �                     @        c       �                    �?R]�M2��?,           0}@       d       �                 ��$:@�=fL�?�            �x@       e       �                    �?�	L �F�?�            `s@        f       }                    �?�<ݚ�?            �F@       g       h                     @:�&���?            �C@        ������������������������       �                     @        i       r                   �7@tk~X��?             B@        j       k                    /@և���X�?             @        ������������������������       �                      @        l       o                    5@���Q��?             @        m       n                 �{@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        p       q                 ���@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        s       t                 ���@\-��p�?             =@        ������������������������       �                     $@        u       |                   �=@���y4F�?             3@       v       {                   �<@������?	             .@       w       z                   @@8�Z$���?             *@       x       y                   @<@z�G�z�?             $@       ������������������������       ��<ݚ�?             "@        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ~                           3@      �?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �@�;���?�            �p@        �       �                     @�J�4�?7            �R@        ������������������������       �                     "@        �       �                 ��@"pc�
�?0            �P@       �       �                 @3�@dP-���?#            �G@        �       �                   �B@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?t��ճC�?!             F@       �       �                 ���@@4և���?             E@        ������������������������       �        	             &@        �       �                    �?��a�n`�?             ?@       �       �                   �<@�t����?             1@       ������������������������       �        	             &@        �       �                    >@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                 ���@@4և���?
             ,@        ������������������������       �                     �?        ������������������������       �        	             *@        ������������������������       �                      @        �       �                    �?D�n�3�?             3@       �       �                   �9@�q�q�?             .@        �       �                   �5@      �?              @       �       �                   �4@      �?             @        ������������������������       �                      @        �       �                 ��L@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �=@և���X�?             @        ������������������������       �                     @        �       �                   @@@      �?             @        �       �                   �?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �9@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                 �?�@�:nR&y�?s            �g@        ������������������������       �                     >@        �       �                   @A@p=
ףp�?a             d@       �       �                    ?@Xny��?I            �^@       �       �                 ���!@�v�\�?=            �Y@        �       �                   �0@4?,R��?             B@        ������������������������       �                     �?        �       �                    �?(N:!���?            �A@       �       �                 pf� @\-��p�?             =@       ������������������������       �                     6@        �       �                   �7@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                     @Pa�	�?*            �P@        �       �                   �(@ 	��p�?             =@        ������������������������       �                     $@        �       �                    �?�KM�]�?             3@       �       �                   �;@      �?             0@       ������������������������       �                     (@        �       �                    =@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                    �B@        �       �                   @@@��Q��?             4@        �       �                    �?r�q��?             @       �       �                 ��i @      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �@@؇���X�?             ,@        ������������������������       �                     @        �       �                    1@z�G�z�?             $@       �       �                 ��%@�q�q�?             @        ������������������������       �                      @        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     C@        �       �                    9@Pi�����?5            �T@        ������������������������       �                      @        �       �                     @l�;�	�?1            �R@       �       �                    �?bKv���?,            @Q@        �       �                    �?     ��?             0@       �       �                   @D@      �?              @       �       �                 ���<@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?Fmq��?!            �J@       �       �                   �>@p�ݯ��?             C@       �       �                 03k:@|��?���?             ;@        ������������������������       �                     @        �       �                   �<@\X��t�?             7@        ������������������������       �                     @        �       �                    R@�E��ӭ�?             2@       �       �                   �J@������?             1@        �       �                   @>@X�<ݚ�?             "@       �       �                   `G@����X�?             @       �       �                   �B@r�q��?             @        ������������������������       �                      @        �       �                   �F@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        �       �                    �?��S���?	             .@       �       �                    D@��
ц��?             *@        �       �                 03�P@؇���X�?             @        ������������������������       �                     @        �       �                   �B@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ���Y@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    >@r�q��?             @       �       �                    ;@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                      @        �                           @���A��?2            �R@                                 2@�Q����?             D@        ������������������������       �        
             ,@                                 �?R�}e�.�?             :@              
                    �?$�q-�?             *@             	                   �?ףp=
�?             $@                               �?@r�q��?             @        ������������������������       �                     @                              �;�p@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                               x�F@��
ц��?
             *@        ������������������������       �                     @                                 @�q�q�?             "@                             ���X@      �?              @                                �?      �?             @        ������������������������       �                     �?                                @F@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?                                 �?ҳ�wY;�?             A@        ������������������������       �                      @                                 �?     ��?             @@        ������������������������       �                     @                                  0@�n_Y�K�?             :@                                 �?�q�q�?             (@                             ���#@���!pc�?             &@        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        !      "                ��T?@؇���X�?
             ,@        ������������������������       �                     @        #      $                   @      �?              @        ������������������������       �                      @        ������������������������       �                     @        �t�bh�h*h-K ��h/��R�(KM%KK��h]�BP       0|@     Pp@      U@      d@      @     �\@       @     �V@             �I@       @      D@              =@       @      &@       @      @       @      @               @       @      �?              �?       @                      @              @      @      7@              &@      @      (@              "@      @      @      @                      @     �S@     �G@     �B@      >@      0@      0@      @              *@      0@      @      (@              @      @       @       @              @       @      �?      �?              �?      �?               @      @               @       @      @               @       @      @       @      �?               @       @      @      @              @      @      @      �?              �?      @                      @      5@      ,@      &@      (@              @      &@      @      &@      @      &@      �?      @      �?       @               @      �?              �?       @              @                       @              @      $@       @      @              @       @      @                       @     �D@      1@      6@      .@              @      6@      &@      2@      $@      *@      @      @              @      @      @      @      @              @      @              �?      @      @      @                      @              �?      @      @      @      �?              �?      @                      @      @      �?      @                      �?      3@       @      *@              @       @               @      @             �v@      Y@     `t@     �P@      q@      B@     �A@      $@      @@      @      @              =@      @      @      @       @               @      @      �?       @      �?                       @      �?      �?              �?      �?              9@      @      $@              .@      @      &@      @      &@       @       @       @      @       @      �?              @                       @      @              @      @              @      @             �m@      :@     �O@      (@      "@              K@      (@     �E@      @       @      �?              �?       @             �D@      @     �C@      @      &@              <@      @      .@       @      &@              @       @               @      @              *@      �?              �?      *@               @              &@       @      $@      @      @      �?      @      �?       @              �?      �?              �?      �?              @              @      @              @      @      �?      �?      �?      �?                      �?       @              �?      @              @      �?              f@      ,@      >@             @b@      ,@      [@      ,@     �W@      @      ?@      @              �?      ?@      @      9@      @      6@              @      @      @                      @      @              P@       @      ;@       @      $@              1@       @      ,@       @      (@               @       @               @       @              @             �B@              *@      @      �?      @      �?      @              @      �?                       @      (@       @      @               @       @      @       @       @               @       @      @              C@              J@      ?@       @              F@      ?@     �E@      :@      &@      @      @      @       @      @       @                      @      �?               @              @@      5@      8@      ,@      *@      ,@              @      *@      $@              @      *@      @      *@      @      @      @      @       @      @      �?       @              @      �?       @      �?      �?                      �?               @       @                      �?      &@               @      @      @      @      �?      @              @      �?      �?      �?                      �?      @              �?      �?      �?                      �?      �?      @      �?      @              �?      �?       @               @     �D@     �@@      3@      5@              ,@      3@      @      (@      �?      "@      �?      @      �?      @               @      �?       @                      �?      @              @              @      @      @              @      @       @      @       @       @              �?       @      �?              �?       @                      @      �?              6@      (@               @      6@      $@      @              0@      $@      @       @      @       @      @                       @      �?              (@       @      @              @       @               @      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�EhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM=huh*h-K ��h/��R�(KM=��h|�B@O         4                   @ ��ʀ_�?�           @�@              =                    �?��W�?�           ��@               0                 pVAH@�ՙ/�?K            �_@                                  �?l��[B��?2            �U@                                  �1@\-��p�?             =@        ������������������������       �                     $@                                   �?���y4F�?             3@        ������������������������       �                     @        	                           �?�	j*D�?             *@       
                        `�@1@      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @                                    @����S��?%             M@                                   (@`�Q��?             9@        ������������������������       �                      @                                   �?��+7��?             7@                                  A@ҳ�wY;�?             1@                               ���<@���Q��?	             .@                               `��,@z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @                                   >@z�G�z�?             @                               03SA@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @               /                    �?���!pc�?            �@@              .                 83�'@�z�G��?             >@               )                   @@�<ݚ�?             ;@       !       "                    5@R���Q�?             4@        ������������������������       �                     @        #       &                 ���@d}h���?             ,@       $       %                   �7@z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        '       (                    9@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        *       +                   �<@և���X�?             @        ������������������������       �                     @        ,       -                    @@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        1       2                    �?$�q-�?            �C@       ������������������������       �                     ;@        3       8                    �?      �?	             (@        4       7                 @�?t@z�G�z�?             @        5       6                   �8@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        9       <                   @C@����X�?             @       :       ;                   �:@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        >       �                     @H\w����?^           ��@        ?       H                   �(@F�����?�            �l@        @       G                    �?@-�_ .�?            �B@       A       B                    @�X�<ݺ?             B@        ������������������������       �                     0@        C       F                   �;@ףp=
�?
             4@        D       E                   �9@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �                     �?        I       �                   �I@�#}���?�            �g@       J       �                    �?@K����?q            �d@       K       \                    :@$/����?U            @`@        L       Q                     �? �o_��?             9@        M       P                 `f�K@z�G�z�?             @        N       O                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        R       U                    �?R���Q�?             4@       S       T                    �?@4և���?
             ,@        ������������������������       �      �?              @        ������������������������       �                     (@        V       W                   �5@�q�q�?             @        ������������������������       �                     �?        X       [                    �?z�G�z�?             @       Y       Z                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ]       �                    �?<W#.m��?C            @Z@       ^       g                    �?���H.�?@             Y@        _       `                     �?�C��2(�?             F@        ������������������������       �                     4@        a       b                   `2@r�q��?             8@       ������������������������       �        	             .@        c       d                    �?X�<ݚ�?             "@        ������������������������       �                     �?        e       f                    <@      �?              @        ������������������������       �                     @        ������������������������       �                     @        h       y                     �?��X��?%             L@       i       p                   �>@�f7�z�?             =@        j       k                 ��$:@�	j*D�?	             *@        ������������������������       �                      @        l       o                   @>@"pc�
�?             &@       m       n                 `f�;@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        q       r                 `fFJ@     ��?             0@       ������������������������       �                     $@        s       t                   @K@      �?             @        ������������������������       �                      @        u       x                    F@      �?             @       v       w                   �@@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        z       �                    ,@�<ݚ�?             ;@       {       |                    @@�	j*D�?	             *@        ������������������������       �                     @        }       ~                 `f�)@���Q��?             $@        ������������������������       �                      @               �                    G@      �?              @       �       �                    C@և���X�?             @       ������������������������       �      �?             @        ������������������������       ��q�q�?             @        ������������������������       �                     �?        �       �                   �7@؇���X�?             ,@        ������������������������       �                     @        �       �                   �:@      �?              @       �       �                    �?�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                 ���[@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?4?,R��?             B@       �       �                    �?���}<S�?             7@       ������������������������       �        
             *@        �       �                    +@z�G�z�?             $@       ������������������������       �                     @        �       �                    A@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                 ���`@�θ�?
             *@       �       �                    �?ףp=
�?             $@       ������������������������       �                      @        �       �                     �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 Ъ�c@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?z�G�z�?             9@        ������������������������       �                     @        �       �                 `fF<@�C��2(�?             6@        ������������������������       �                     (@        �       �                     �?z�G�z�?             $@       �       �                    �?�<ݚ�?             "@       �       �                   @>@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    /@��O��?�            �s@        �       �                    �?ףp=
�?             $@        ������������������������       �                     @        �       �                 033<@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       +                  @@@�=A�F�?�             s@       �                         �>@����F��?�            �m@       �       �                 �1@�θ�?�            �k@        �       �                    �?�Z4���?.            �P@       �       �                 �@��~R���?,            �O@        �       �                    �?���Q��?             .@        ������������������������       �                     @        �       �                    �?�eP*L��?	             &@        ������������������������       �                     �?        �       �                    7@      �?             $@        ������������������������       �                     @        �       �                 ���@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�q�q�?!             H@        �       �                    �?b�2�tk�?             2@       �       �                   �5@�	j*D�?	             *@        �       �                  s�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                  ��@z�G�z�?             $@        ������������������������       �                     �?        �       �                    �?�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        �       �                 ���@���Q��?             @        ������������������������       �                     �?        �       �                    4@      �?             @        ������������������������       �                      @        �       �                   �7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �<@ףp=
�?             >@       �       �                   �;@ 	��p�?             =@       �       �                 �?$@؇���X�?
             ,@       ������������������������       �                     &@        �       �                   �6@�q�q�?             @        ������������������������       �                     �?        �       �                   �9@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             .@        ������������������������       �                     �?        �       �                   �7@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �                          �?z���=��?a            @c@       �                       �T)D@�MI8d�?]            �b@       �       �                    �?`	�<��?[            �a@        �       �                    �?X�Cc�?             <@        �       �                 03�'@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?`�Q��?             9@       �       �                    �?���N8�?             5@       �       �                    �?z�G�z�?             .@       �       �                 ��&@ףp=
�?	             $@       ������������������������       �                     "@        ������������������������       �                     �?        �       �                 �̬)@���Q��?             @        ������������������������       �                      @        �       �                    9@�q�q�?             @        ������������������������       �                     �?        �       �                    ;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �;@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 �?�@4�0_���?C            @\@        ������������������������       �                     ?@        �                          �?�<p���?0            �T@       �       �                    �?H%u��?,            �R@        ������������������������       �                     $@        �                         �:@��ɉ�?'            @P@        �                          �? 	��p�?             =@       �                       ��Y @h�����?             <@                               @3�@�C��2(�?             &@        ������������������������       �                     �?                                �3@ףp=
�?             $@                                �1@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �        
             1@        ������������������������       �                     �?        	                         �?tk~X��?             B@       
                      ��) @�'�`d�?            �@@        ������������������������       �                     ,@                              ��)"@p�ݯ��?
             3@                              pf� @r�q��?             @        ������������������������       �                      @                                �;@      �?             @        ������������������������       �                     @        ������������������������       �                     �?                                 (@8�Z$���?             *@                               �<@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �����X�?             @                                 �?�q�q�?             @                                �?      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @              *                   �?b�2�tk�?	             2@              !                �?�@ҳ�wY;�?             1@        ������������������������       �                     @        "      )                `��(@�eP*L��?             &@       #      $                   �?      �?              @        ������������������������       �                     �?        %      &                  �?@����X�?             @        ������������������������       �                      @        '      (                @3�@���Q��?             @       ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ,      3                @3�@��ɉ�?+            @P@        -      .                �?�@��S�ۿ?             >@       ������������������������       �                     8@        /      2                  �D@�q�q�?             @       0      1                   C@z�G�z�?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                    �A@        5      6                ��	5@t��ճC�?             F@        ������������������������       �                      @        7      <                   @�Ń��̧?             E@        8      9                   @؇���X�?             @       ������������������������       �                     @        :      ;                ���A@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                    �A@        �t�b�      h�h*h-K ��h/��R�(KM=KK��h]�B�       �|@     �o@     z@     `o@      H@     �S@     �F@      E@      @      9@              $@      @      .@              @      @      "@      @      @      @                      @              @     �D@      1@      1@       @               @      1@      @      &@      @      "@      @       @       @               @       @              �?      @      �?       @               @      �?                       @       @              @              8@      "@      5@      "@      5@      @      1@      @      @              &@      @       @       @               @       @              @      �?      �?               @      �?      @      @      @              �?      @              @      �?                      @      @              @      B@              ;@      @      "@      �?      @      �?      �?      �?                      �?              @       @      @       @       @               @       @                      @     w@     �e@      _@      Z@     �A@       @      A@       @      0@              2@       @       @       @       @                       @      $@              �?             @V@     �Y@     @Q@     @X@      P@     �P@      2@      @      �?      @      �?      �?              �?      �?                      @      1@      @      *@      �?      �?      �?      (@              @       @              �?      @      �?       @      �?              �?       @               @              G@     �M@      E@      M@      @      D@              4@      @      4@              .@      @      @              �?      @      @      @                      @      C@      2@      1@      (@      @      "@       @               @      "@       @      @              @       @                      @      *@      @      $@              @      @               @      @      �?      �?      �?      �?                      �?       @              5@      @      "@      @      @              @      @       @              @      @      @      @       @       @      �?       @      �?              (@       @      @              @       @      @       @      @                       @       @              @      �?      @                      �?      @      ?@       @      5@              *@       @       @              @       @      �?       @                      �?      @      $@      �?      "@               @      �?      �?              �?      �?               @      �?       @                      �?      4@      @              @      4@       @      (@               @       @      @       @      @       @               @      @              @              �?             �n@     @Q@      �?      "@              @      �?      @              @      �?             �n@      N@     �f@      M@     @e@     �I@      E@      9@      D@      7@      @      "@              @      @      @      �?              @      @      @               @      @              @       @              A@      ,@      @      &@      @      "@       @      �?              �?       @               @       @      �?              �?       @               @      �?              @       @              �?      @      �?       @              �?      �?              �?      �?              ;@      @      ;@       @      (@       @      &@              �?       @              �?      �?      �?      �?                      �?      .@                      �?       @       @       @                       @      `@      :@      _@      8@     �^@      3@      2@      $@      �?       @      �?                       @      1@       @      0@      @      (@      @      "@      �?      "@                      �?      @       @       @              �?       @              �?      �?      �?      �?                      �?      @       @               @      @              �?      @              @      �?              Z@      "@      ?@             @R@      "@     �P@      "@      $@              L@      "@      ;@       @      ;@      �?      $@      �?      �?              "@      �?       @      �?      �?              �?      �?      @              1@                      �?      =@      @      :@      @      ,@              (@      @      �?      @               @      �?      @              @      �?              &@       @      @       @      @                       @      @              @              @               @      @      @       @       @       @               @       @               @              &@      @      &@      @      @              @      @       @      @              �?       @      @               @       @      @       @      �?               @      @                      �?     �O@       @      <@       @      8@              @       @      @      �?       @               @      �?              �?     �A@             �D@      @               @     �D@      �?      @      �?      @              �?      �?              �?      �?             �A@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ4�phG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B�A         h                     @@?�p�?�           @�@               A                 03�I@(�ruX��?�            0s@                                  �?���_�?v            @g@                                   �?@3����?)             K@        ������������������������       �                     *@                                   �?��Y��]�?!            �D@                                 �9@ ��WV�?             :@                                  �3@r�q��?             @       	       
                   �6@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     4@        ������������������������       �                     .@               8                    �?�������?M            �`@              )                     �? ��(��?B            @\@                                ��I*@�J��%�?            �H@        ������������������������       �                      @                                03k:@hP�vCu�?            �D@        ������������������������       �                     @               (                    R@<ݚ)�?             B@              !                    �?r�q��?             >@                                   �L@�<ݚ�?             "@                                 �E@����X�?             @                                  =@r�q��?             @                               �ܵ<@�q�q�?             @        ������������������������       �                     �?                                03SA@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        "       '                   �<@؇���X�?             5@        #       &                 ��yC@�q�q�?             "@       $       %                 `fF<@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     (@        ������������������������       �                     @        *       1                    �?      �?'             P@       +       ,                    �? qP��B�?            �E@        ������������������������       �                     @        -       0                    &@P�Lt�<�?             C@        .       /                   �H@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     =@        2       7                    @@؇���X�?	             5@        3       4                   �7@և���X�?             @        ������������������������       �                     �?        5       6                   �<@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     ,@        9       >                 �DpB@p�ݯ��?             3@       :       ;                     �?8�Z$���?             *@        ������������������������       �                     �?        <       =                    +@r�q��?             (@        ������������������������       �                      @        ������������������������       �                     $@        ?       @                   �>@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        B       g                    O@�#DwKd�?G            @^@       C       D                    �?�θ�?E            @]@       ������������������������       �        (            �Q@        E       F                   �1@�[�IJ�?            �G@        ������������������������       �                     "@        G       N                    �?p9W��S�?             C@        H       M                   �;@�r����?             .@       I       L                 Ј@S@����X�?             @        J       K                     �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        O       d                    �?�û��|�?             7@       P       c                     �?��Q��?             4@       Q       X                   �;@p�ݯ��?             3@        R       W                 �U�X@���Q��?             @       S       V                 0�"K@      �?             @        T       U                    7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        Y       ^                   �G@����X�?	             ,@       Z       ]                 03�M@�����H�?             "@        [       \                   @K@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        _       `                   �H@���Q��?             @        ������������������������       �                      @        a       b                 `f^@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        e       f                     @�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        i       �                    �?���iz�?�            Py@        j       {                    �?Υf���?D            �^@        k       r                   �6@�	j*D�?            �C@        l       q                    0@�G�z��?	             4@       m       n                    �?ףp=
�?             $@       ������������������������       �                     @        o       p                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        s       t                    :@�}�+r��?             3@        ������������������������       �                      @        u       z                    �?�IєX�?             1@        v       y                    �?      �?              @        w       x                 �%@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        |       �                    �?F~��7�?/            �T@        }       �                    @<=�,S��?            �A@       ~       �                   �;@�q�q�?            �@@              �                    �?��+7��?             7@       �       �                    9@     ��?             0@       �       �                    �?      �?             $@       �       �                 �[$@      �?              @       �       �                 P��@�q�q�?             @        ������������������������       �                     �?        �       �                 @�"@���Q��?             @       �       �                  � @      �?             @       �       �                    4@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �&@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                 `f7@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �>@      �?             $@       �       �                    =@����X�?             @        ������������������������       �                     �?        �       �                 @3#%@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                    @r�qG�?             H@       �       �                    �?�^�����?            �E@       �       �                    �?d��0u��?             >@       �       �                    @���Q��?
             4@       �       �                 �̬)@�t����?	             1@        ������������������������       �                     @        �       �                 ��1@�n_Y�K�?             *@       �       �                 @3�/@X�<ݚ�?             "@        ������������������������       �                     �?        �       �                    ;@      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                     @�z�G��?             $@       �       �                 `f�.@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                 ���1@8�Z$���?             *@        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �                     @        �       �                    �?P�I;l�?�            �q@        �       �                    5@:ɨ��?            �@@        �       �                 �{@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   @@8�Z$���?             :@       �       �                   �7@��s����?             5@        �       �                 ���@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                 ���@      �?             0@       ������������������������       �                     "@        �       �                   @<@����X�?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @ĭ����?�            @o@        �       �                    @�q�q�?             (@       �       �                    @����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �<@T�W2��?�            �m@       �       �                  ��	@�YX�Z�?e            �d@        ������������������������       �                     �?        �       �                    �?x�}���?d            �d@       �       �                    �?���7�?]            @c@       �       �                    ;@`�q�0ܴ?U            �a@       �       �                    �?�F��O�?+            @R@       �       �                 `�B@�8��8��?*             R@       �       �                 ���@ >�֕�?)            �Q@        �       �                    �?z�G�z�?             $@       �       �                 �&b@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?(;L]n�?#             N@       �       �                 �1@@3����?              K@        �       �                 �?$@�8��8��?	             (@       ������������������������       �                     $@        �       �                   �5@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     E@        �       �                    5@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        *             Q@        �       �                 ���2@$�q-�?             *@        �       �                 xFT$@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     (@        �                          @@@�ӖF2��?+            �Q@        �       �                   �=@�G��l��?             5@        �       �                    �?���Q��?             @        ������������������������       �                      @        �       �                 ���"@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �?@     ��?             0@        ������������������������       �                      @        �       �                 �!B@      �?
             ,@       �       �                 �Y5@���|���?             &@        ������������������������       �                      @        �       �                 pf�'@X�<ݚ�?             "@       �       �                 @3�@և���X�?             @       �       �                   �@���Q��?             @        ������������������������       �                     �?        �       �                 �?�@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @                                �E@p���?             I@       ������������������������       �                     ?@                              P�@�}�+r��?	             3@       ������������������������       �                     (@                                �G@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h*h-K ��h/��R�(KMKK��h]�Bp       �{@     �p@      a@     @e@     �Z@      T@      �?     �J@              *@      �?      D@      �?      9@      �?      @      �?       @              �?      �?      �?              @              4@              .@     @Z@      ;@     @W@      4@     �@@      0@       @              9@      0@              @      9@      &@      9@      @      @       @      @       @      @      �?       @      �?      �?              �?      �?              �?      �?              @                      �?       @              2@      @      @      @      �?      @      �?                      @      @              (@                      @      N@      @      E@      �?      @             �B@      �?       @      �?       @                      �?      =@              2@      @      @      @      �?              @      @      @                      @      ,@              (@      @      &@       @      �?              $@       @               @      $@              �?      @              @      �?              ?@     �V@      ;@     �V@             �Q@      ;@      4@              "@      ;@      &@      *@       @      @       @       @       @               @       @              @               @              ,@      "@      *@      @      (@      @       @      @      �?      @      �?      �?      �?                      �?               @      �?              $@      @       @      �?      �?      �?      �?                      �?      @               @      @               @       @      �?       @                      �?      �?              �?       @               @      �?              @             0s@     �X@      N@      O@      (@      ;@      &@      "@      �?      "@              @      �?       @      �?                       @      $@              �?      2@               @      �?      0@      �?      @      �?      �?              �?      �?                      @              "@      H@     �A@      *@      6@      &@      6@      @      1@      @      &@      @      @      @      @       @      @              �?       @      @       @       @      �?       @      �?                       @      �?                      �?       @              �?      �?      �?                      �?              @      �?      @              @      �?              @      @      @       @      �?              @       @      @                       @              @       @             �A@      *@      >@      *@      3@      &@      (@       @      (@      @      @               @      @      @      @              �?      @      @      @                      @      @                      @      @      @       @      @       @                      @      @              &@       @               @      &@              @             �n@      B@      7@      $@      �?      @      �?                      @      6@      @      1@      @      @       @               @      @              ,@       @      "@              @       @      @       @      �?              @              l@      :@      @      @      @       @               @      @                      @     `k@      3@     �c@       @              �?     �c@      @     `b@      @     �`@      @     �P@      @     �P@      @     �P@      @       @       @      @       @      @                       @      @              M@       @     �J@      �?      &@      �?      $@              �?      �?              �?      �?              E@              @      �?              �?      @                       @      �?              Q@              (@      �?       @      �?       @                      �?      $@              (@              N@      &@      &@      $@       @      @               @       @      �?       @                      �?      "@      @       @              @      @      @      @       @              @      @      @      @      @       @              �?      @      �?      �?               @      �?               @       @                      @     �H@      �?      ?@              2@      �?      (@              @      �?              �?      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJLxhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM7huh*h-K ��h/��R�(KM7��h|�B�M         >                    �?^IB�A��?�           @�@               %                     @r���@�?J            �Z@              
                   �;@:-�.A�?+            �P@               	                    �?���}<S�?             7@                                  �?�r����?
             .@        ������������������������       �                     @                                 ��^@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @                                p�H@�zv�X�?             F@                                   �?     ��?
             0@        ������������������������       �                     �?                                    �?������?	             .@       ������������������������       �                     @                                   �?X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @                                    �?d}h���?             <@                                  �?��<b���?             7@       ������������������������       �                     (@                                 �}S@�eP*L��?             &@        ������������������������       �                      @                                   �?X�<ݚ�?             "@                                 �?@�q�q�?             @        ������������������������       �                      @                                �;|r@      �?             @        ������������������������       �                      @        ������������������������       �                      @                                  �H@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        !       $                    �?z�G�z�?             @       "       #                   �E@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        &       7                 033.@�G�z��?             D@       '       ,                    �?8^s]e�?             =@        (       +                    7@���Q��?             $@       )       *                 P��+@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        -       .                   @@�S����?             3@       ������������������������       �        	             (@        /       6                    ?@և���X�?             @       0       5                   �<@���Q��?             @       1       2                 83##@�q�q�?             @        ������������������������       �                     �?        3       4                    4@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        8       =                    �?"pc�
�?	             &@        9       <                    �?�q�q�?             @       :       ;                   �2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ?                          �?��\��?z           �@       @       �                 0#�9@�����?            �|@       A       h                     @dd��G��?�            �u@        B       C                     �?�ucQ?-�?8            @U@        ������������������������       �                     @        D       G                    �?�q�q�?4            �S@        E       F                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        H       M                    �?`�Q��?1            �R@        I       J                   �'@�X�<ݺ?             2@        ������������������������       �                     @        K       L                    :@�C��2(�?	             &@        ������������������������       ��q�q�?             @        ������������������������       �                      @        N       e                    M@���5��?#            �L@       O       d                    �?lGts��?!            �K@       P       Q                    @�q��/��?            �H@        ������������������������       �                     @        R       c                   @F@��2(&�?             F@       S       b                    C@b�h�d.�?            �A@       T       Y                    &@      �?             @@        U       X                   �5@"pc�
�?             &@        V       W                   �1@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        Z       [                   �;@�����?             5@        ������������������������       �                     (@        \       ]                 `fF)@�<ݚ�?             "@        ������������������������       �                     �?        ^       a                   �*@      �?              @       _       `                    =@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     "@        ������������������������       �                     @        f       g                   �P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        i       �                    �? 0|zJ�?�            Pp@        j       q                  ��@     ��?             H@        k       p                 @3�@r�q��?             @       l       m                   �8@�q�q�?             @        ������������������������       �                     �?        n       o                 ���@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        r                           �?�G��l��?             E@       s       ~                   �>@�5��?             ;@       t       }                 pF @r�q��?             8@       u       x                    �?      �?             6@        v       w                   �5@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        y       |                 ��(@r�q��?	             (@       z       {                   �<@"pc�
�?             &@       ������������������������       �ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                 03�7@���Q��?             .@       �       �                    �?X�Cc�?             ,@       ������������������������       �                     "@        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�OJ�+�?�            �j@       �       �                    O@��vA��?�            `i@       �       �                    �?T�{J�~�?�            @i@        �       �                    3@J�8���?             =@        ������������������������       �                      @        �       �                   �7@l��
I��?             ;@        �       �                 pf&@�q�q�?             (@        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?z�G�z�?	             .@        ������������������������       �                     @        �       �                 @3S)@      �?              @        ������������������������       �                     @        �       �                   �=@      �?             @        ������������������������       �                      @        �       �                   �@@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 �1@�߄��?m            �e@        �       �                 �?$@&y�X���?&             M@       �       �                 @3�@ i���t�?"            �H@        �       �                   �>@�q�q�?             @        �       �                    6@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?Du9iH��?            �E@       �       �                   �>@�˹�m��?             C@       �       �                    7@�LQ�1	�?             7@        ������������������������       �        	             "@        �       �                   �8@d}h���?	             ,@        ������������������������       �                     �?        �       �                    ;@8�Z$���?             *@        ������������������������       �                     @        �       �                 pf�@z�G�z�?             $@       ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �        	             .@        ������������������������       �                     @        �       �                   �;@�q�q�?             "@       �       �                   �5@؇���X�?             @        ������������������������       �                     @        �       �                   �8@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                 �?�@������?G            �\@        �       �                    ?@������?             B@       ������������������������       �                     ?@        �       �                   �@z�G�z�?             @        �       �                    D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                 @3�@p#�����?2            �S@        �       �                    :@      �?             $@        ������������������������       �                     �?        �       �                   �?@X�<ݚ�?             "@        ������������������������       �                     �?        �       �                   �A@      �?              @        ������������������������       �      �?              @        ������������������������       �      �?             @        �       �                 ��) @���}<S�?,            @Q@        �       �                    ?@XB���?             =@       ������������������������       �                     5@        �       �                   �@@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ��y @      �?             D@        ������������������������       �                      @        �       �                    �?�˹�m��?             C@       �       �                    (@�#-���?            �A@       �       �                   �8@ףp=
�?             >@        ������������������������       �                     *@        �       �                 ���"@@�0�!��?	             1@       �       �                 ���!@�r����?             .@       �       �                   �;@r�q��?             (@        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �                     @        �       �                    ?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        �       �                    �?�X���?D             \@        ������������������������       �                     I@        �       �                     @�&�5y�?*             O@       �       �                   @J@4և����?%             L@       �       �                    �?�7����?            �G@       �       �                   @H@�q�q�?             8@       �       �                 `f�;@��+7��?             7@       �       �                   �F@��
ц��?             *@       �       �                 ��$:@�eP*L��?             &@        ������������������������       �                      @        �       �                   �A@�q�q�?             "@        ������������������������       ����Q��?             @        �       �                   �E@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �                     �?        �       �                    H@��+7��?             7@       �       �                    �?�GN�z�?             6@       �       �                    D@      �?             4@       �       �                     �?�q�q�?	             .@       �       �                   �B@�q�q�?             (@       �       �                 `f�N@���|���?             &@       �       �                 `fFJ@և���X�?             @        ������������������������       �                      @        �       �                    7@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@                                  ;@�q�q�?             @        ������������������������       �                      @                                 >@      �?             @        ������������������������       �                      @        ������������������������       �                      @              (                  �9@��7���?Z            `b@                             03�;@4�	~���?.            @Q@                               �0@�p ��?            �D@                                @�θ�?             :@       	                         �?ףp=
�?             4@       
                          @      �?
             0@        ������������������������       �                     "@                                 @����X�?             @                                �?      �?             @        ������������������������       �                     �?                              pf�0@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @                                 �?�q�q�?             @        ������������������������       �                     @                              032@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     .@                              ��T?@և���X�?             <@        ������������������������       �                      @                                 �?���Q��?             4@        ������������������������       �                     @              %                     @��S���?             .@              "                    @      �?              @               !                   �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        #      $                   5@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        &      '                   @և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        )      6                03�X@�q�q�?,            �S@       *      +                ��,2@������?'             Q@        ������������������������       �                     $@        ,      1                   �?�c�Α�?!             M@       -      .                    @      �?             >@        ������������������������       �                     &@        /      0                ���4@���y4F�?	             3@        ������������������������       �                     @        ������������������������       �                     .@        2      3                  `B@h�����?             <@       ������������������������       �                     6@        4      5                   C@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        �t�bh�h*h-K ��h/��R�(KM7KK��h]�Bp       �z@     �q@     �D@     �P@      3@      H@       @      5@       @      *@              @       @      @              @       @                       @      1@      ;@      &@      @              �?      &@      @      @              @      @              @      @              @      6@      @      2@              (@      @      @               @      @      @      @       @       @               @       @       @                       @      �?       @               @      �?              �?      @      �?      �?              �?      �?                      @      6@      2@      4@      "@      @      @      @       @               @      @                      @      0@      @      (@              @      @       @      @       @      �?      �?              �?      �?              �?      �?                       @       @               @      "@       @      �?      �?      �?      �?                      �?      �?                       @      x@     �k@     `s@     �b@     �p@     @T@     �M@      :@      @              J@      :@      �?       @               @      �?             �I@      8@      �?      1@              @      �?      $@      �?       @               @      I@      @     �H@      @     �E@      @      @              C@      @      =@      @      <@      @      "@       @      �?       @      �?                       @       @              3@       @      (@              @       @      �?              @       @      @       @               @      @              �?              �?       @      "@              @              �?      �?              �?      �?             �i@     �K@      ;@      5@      @      �?       @      �?      �?              �?      �?      �?                      �?      @              6@      4@      0@      &@      *@      &@      &@      &@      �?      "@      �?                      "@      $@       @      "@       @      "@      �?              �?      �?               @              @              @      "@      @      "@              "@      @              �?             `f@      A@      e@      A@      e@     �@@      3@      $@               @      3@       @      @      @              @      @              (@      @      @              @      @      @              �?      @               @      �?      �?      �?                      �?     �b@      7@     �G@      &@      F@      @      @       @      �?       @      �?                       @      @              D@      @     �A@      @      4@      @      "@              &@      @              �?      &@       @      @               @       @      @              �?       @      .@              @              @      @      �?      @              @      �?      @      �?                      @       @             �Y@      (@     �A@      �?      ?@              @      �?      �?      �?              �?      �?              @              Q@      &@      @      @      �?              @      @              �?      @      @      �?      �?      @      @     �O@      @      <@      �?      5@              @      �?              �?      @             �A@      @               @     �A@      @      @@      @      ;@      @      *@              ,@      @      *@       @      $@       @               @      $@              @              �?      �?              �?      �?              @              @                      �?      $@             �F@     �P@              I@     �F@      1@     �E@      *@      A@      *@      1@      @      1@      @      @      @      @      @       @              @      @       @      @      �?      @              �?      �?       @       @              $@                      �?      1@      @      1@      @      .@      @      $@      @      @      @      @      @      @      @       @              �?      @      �?                      @      @                      �?      @              @               @                      �?      "@               @      @               @       @       @       @                       @     �R@     @R@      6@     �G@      @     �A@      @      4@       @      2@       @      ,@              "@       @      @       @       @              �?       @      �?              �?       @                      @              @      @       @      @              �?       @               @      �?                      .@      0@      (@       @               @      (@              @       @      @      @      @       @      �?       @                      �?       @      @       @                      @      @      @              @      @              J@      :@      J@      0@      $@              E@      0@      .@      .@              &@      .@      @              @      .@              ;@      �?      6@              @      �?              �?      @                      $@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJW��8hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM9huh*h-K ��h/��R�(KM9��h|�B@N         j                    �?��!h
��?�           @�@                                    @Ȩ�I��?�            �p@                                  �? 7���B�?Q            �`@                                 �;@ rpa�?7            @W@               
                   �9@r�q��?             8@              	                 ��*@�C��2(�?             6@                                  �'@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        
             3@        ������������������������       �                      @                                   �?@	tbA@�?*            @Q@                                  �?��Y��]�?            �D@                                  �G@ףp=
�?             $@       ������������������������       �                     @                                ,w�U@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     ?@        ������������������������       �                     <@        ������������������������       �                     E@               c                 ��Y7@      �?L            @`@                               ���@�5��?@             [@                                 �[@�8��8��?	             (@       ������������������������       �                     @                                  �8@z�G�z�?             @        ������������������������       �                      @                                 ��@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @               6                    �?r�q��?7             X@                /                    �?     ��?             @@       !       &                   �5@�q�q�?             ;@        "       #                    �?      �?              @        ������������������������       �                     @        $       %                    2@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        '       .                 03�'@�S����?
             3@       (       -                 pF @�θ�?             *@       )       *                    9@r�q��?             (@        ������������������������       �                     �?        +       ,                 �&B@"pc�
�?             &@       ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        0       5                    �?���Q��?             @       1       4                   �<@      �?             @       2       3                    -@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        7       V                 `f�%@      �?%             P@       8       U                    �?���Q��?             D@       9       T                 �[$@�'�=z��?            �@@       :       S                    �?П[;U��?             =@       ;       R                  �m#@���>4��?             <@       <       =                 ��@r�q��?             8@        ������������������������       �                      @        >       O                 `��!@      �?             6@       ?       H                 �?�@     ��?
             0@        @       C                 �&B@X�<ݚ�?             "@        A       B                   �7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        D       G                   �@�q�q�?             @       E       F                    4@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        I       J                   �8@����X�?             @        ������������������������       �                     �?        K       L                 @3�@r�q��?             @        ������������������������       �                     @        M       N                 ��� @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        P       Q                    I@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        W       b                 ���4@�q�q�?             8@       X       a                    �?���N8�?             5@        Y       Z                    5@X�<ݚ�?             "@        ������������������������       �                     @        [       \                 ��Y.@�q�q�?             @        ������������������������       �                     �?        ]       ^                 @3�/@z�G�z�?             @        ������������������������       �                     �?        _       `                    ;@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        ������������������������       �                     @        d       e                    @���7�?             6@       ������������������������       �        	             1@        f       i                    @z�G�z�?             @       g       h                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        k       �                    �?>���_�?           �{@        l       w                   @@�sly47�?+            �R@        m       v                    �?؇���X�?             5@       n       q                    8@r�q��?             2@        o       p                 �{@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        r       u                   `B@��S�ۿ?	             .@       s       t                 ���@$�q-�?             *@        ������������������������       �                     @        ������������������������       �ףp=
�?             $@        ������������������������       �                      @        ������������������������       �                     @        x       y                   �6@��}*_��?             K@        ������������������������       �                     @        z       �                  I>@�7����?            �G@        {       �                    �?R���Q�?             4@       |       �                 ���4@�z�G��?             $@       }       �                 pf�&@      �?              @       ~       �                    ?@����X�?             @              �                   �<@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        �       �                 �D�@@��}*_��?             ;@        ������������������������       �                     @        �       �                 xCQ@��+7��?             7@        ������������������������       �                      @        �       �                  �}S@���Q��?	             .@        ������������������������       �                      @        �       �                 p�w@�	j*D�?             *@       �       �                    �?      �?             (@        ������������������������       �                     @        �       �                 ��+T@���Q��?             @        ������������������������       �                      @        �       �                   �U@�q�q�?             @        ������������������������       �                     �?        �       �                 ��>Y@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ��l1@����;�?�            @w@       �       �                 �?�@P��4���?�            �o@        �       �                    �?��	,UP�?A             W@        �       �                  s�@      �?             0@       ������������������������       �                     "@        �       �                   �=@؇���X�?             @       ������������������������       �      �?             @        ������������������������       �                     @        �       �                    �?�}�+r��?6             S@       �       �                   �;@0z�(>��?3            �Q@        �       �                   �:@�LQ�1	�?             7@       �       �                 @33@���N8�?             5@        ������������������������       �                     �?        ������������������������       �                     4@        ������������������������       �                      @        ������������������������       �        !             H@        �       �                    5@z�G�z�?             @        ������������������������       �                     @        �       �                 �&B@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 @3�@B�xX�?`            `d@        �       �                    �?      �?             0@       �       �                   �4@և���X�?
             ,@        ������������������������       �                     �?        �       �                   �D@�n_Y�K�?	             *@       �       �                    :@�q�q�?             (@        ������������������������       �                      @        �       �                   �?@���Q��?             $@        ������������������������       �                     �?        �       �                   �A@�q�q�?             "@       ������������������������       ����Q��?             @        ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�q��/��?U            `b@        ������������������������       �                     @        �       �                   �*@������?R            �a@       �       �                    $@�SM:$�?C            @\@        ������������������������       �                     �?        �       �                    �?>4և�z�?B             \@       �       �                    �?��#:���?A            �[@       �       �                 ���"@BMĹ��??             [@       �       �                 ��i @lGts��?             �K@       �       �                   �4@(L���?            �E@        �       �                   �1@���|���?             &@        ������������������������       �      �?              @        ������������������������       ��q�q�?             @        �       �                    ?@      �?             @@       ������������������������       �                     9@        �       �                   �@@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     (@        �       �                     @ {��e�?            �J@       �       �                   �;@t/*�?            �G@        �       �                    5@���}<S�?             7@        �       �                    &@z�G�z�?             $@        �       �                   �1@�q�q�?             @        ������������������������       �                      @        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     *@        �       �                 `f�)@      �?             8@        �       �                   @L@r�q��?             @       ������������������������       �                     @        �       �                   �P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    =@�E��ӭ�?	             2@        ������������������������       �                      @        �       �                    G@     ��?             0@       �       �                   @D@���!pc�?             &@       �       �                    @@      �?              @        ������������������������       �                      @        �       �                   @B@r�q��?             @       ������������������������       �      �?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                     @        �       �                   �:@      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     ;@        �       "                   �?2�ަ��?M            @]@       �                           @L�w�=�?,            �Q@       �       �                 ��$:@����S��?&             M@        �       �                   �@@@4և���?             ,@        �       �                   �>@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        �       �                    �?���|���?             F@        ������������������������       �                     �?        �                          �?�lg����?            �E@       �                         �J@      �?             8@       �       
                   H@���Q��?             4@       �       	                  �F@X�<ݚ�?             2@       �       �                 03k:@j���� �?
             1@        ������������������������       �                      @        �                         �A@��S���?             .@       �                         @@@���Q��?             $@       �                       `fF<@      �?              @                                @B@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @                                �<@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @                                �E@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                 D@���y4F�?
             3@                                �?�q�q�?             (@                             `fFJ@���Q��?             $@        ������������������������       �                      @                                 >@      �?              @                                <@z�G�z�?             @                                7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @              !                  �A@      �?             (@                                 �?���Q��?             $@                             �T)D@և���X�?             @        ������������������������       �                     @                                 >@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        #      2                   @�*/�8V�?!            �G@       $      %                   $@�5��?             ;@        ������������������������       �                     @        &      -                   �?z�G�z�?             4@       '      ,                   D@�r����?
             .@        (      +                    �?����X�?             @        )      *                   �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        .      1                   @���Q��?             @       /      0                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        3      8                   @P���Q�?             4@        4      7                ���A@r�q��?             @        5      6                ��A>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             ,@        �t�b� %     h�h*h-K ��h/��R�(KM9KK��h]�B�       �z@     �q@     �Q@     `h@      @     @`@      @      V@      @      4@       @      4@       @      �?              �?       @                      3@       @              �?      Q@      �?      D@      �?      "@              @      �?       @      �?                       @              ?@              <@              E@     @P@     @P@      F@      P@      �?      &@              @      �?      @               @      �?       @      �?                       @     �E@     �J@      &@      5@      "@      2@      @       @      @              �?       @               @      �?              @      0@      @      $@       @      $@              �?       @      "@       @      @              @      �?                      @       @      @      �?      @      �?      �?              �?      �?                       @      �?              @@      @@      8@      0@      1@      0@      *@      0@      *@      .@      *@      &@       @              &@      &@      @      "@      @      @      �?       @               @      �?              @       @      @       @      @                       @      �?               @      @      �?              �?      @              @      �?      �?      �?                      �?      @       @      @                       @              @              �?      @              @               @      0@      @      0@      @      @      @               @      @      �?              �?      @              �?      �?      @      �?                      @              (@      @              5@      �?      1@              @      �?      �?      �?              �?      �?              @             �v@     �U@      J@      7@      2@      @      .@      @      �?       @      �?                       @      ,@      �?      (@      �?      @              "@      �?       @              @              A@      4@              @      A@      *@      1@      @      @      @      @      @      @       @       @       @       @                       @      @                      �?       @              $@              1@      $@              @      1@      @       @              "@      @               @      "@      @      "@      @      @               @      @               @       @      �?      �?              �?      �?              �?      �?                      �?     @s@      P@     @l@      =@     �U@      @      .@      �?      "@              @      �?      @      �?      @              R@      @      Q@      @      4@      @      4@      �?              �?      4@                       @      H@              @      �?      @              �?      �?              �?      �?             `a@      8@      $@      @       @      @              �?       @      @       @      @       @              @      @              �?      @      @      @       @      @      �?              �?       @              `@      2@      @             �^@      2@     �W@      2@              �?     �W@      1@     @W@      1@     �V@      1@     �H@      @     �B@      @      @      @      @      @       @      �?      >@       @      9@              @       @               @      @              (@              E@      &@     �C@       @      5@       @       @       @      @       @       @               @       @      @              *@              2@      @      @      �?      @              �?      �?              �?      �?              *@      @               @      *@      @       @      @      @      �?       @              @      �?      @      �?       @              �?       @      @              @      @      @                      @       @               @              ;@             �T@     �A@     �G@      7@     �D@      1@      *@      �?      @      �?      @                      �?      $@              <@      0@      �?              ;@      0@      (@      (@       @      (@       @      $@      @      $@               @      @       @      @      @      @      @       @       @      �?              �?       @       @       @               @       @               @              �?      @              @      �?              �?                       @      @              .@      @       @      @      @      @       @              @      @      @      �?      �?      �?      �?                      �?      @                      @       @              @              @      @      @      @      @      @      @              �?      @      �?                      @              @       @             �A@      (@      0@      &@              @      0@      @      *@       @      @       @      �?       @      �?                       @      @               @              @       @       @       @               @       @              �?              3@      �?      @      �?      �?      �?      �?                      �?      @              ,@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ��UhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM/huh*h-K ��h/��R�(KM/��h|�B�K         h                    �?����?�           @�@                                   )@��PN���?�             l@                                   �?��
ц��?             :@        ������������������������       �                     @                                03�<@���|���?             6@                                   @��
ц��?	             *@                                 �&@�z�G��?             $@        ������������������������       �                     �?        	       
                    �?�<ݚ�?             "@        ������������������������       �                     @                                `f7@���Q��?             @        ������������������������       �                      @                                   !@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                   �?�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @               g                    @�<;P�?�            �h@              d                 p�H@8�v�l�?~             h@              c                    J@�E��ӭ�?S            �_@                               ���@*AA,�P�?P            @^@        ������������������������       �                     *@               &                     @�Sb(�	�?H             [@                                   �?�C��2(�?             F@                                0Cd=@      �?             @                                ��@5@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @                !                    �?P�Lt�<�?             C@       ������������������������       �                     :@        "       %                   �7@�8��8��?             (@        #       $                   �<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        '       >                    �?     ��?+             P@        (       -                   �6@�	j*D�?             :@        )       ,                 �{&@      �?             @        *       +                 @�@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        .       =                   �<@�GN�z�?             6@       /       8                    �?�d�����?             3@        0       1                    �?�q�q�?             "@        ������������������������       �                      @        2       3                    �?؇���X�?             @        ������������������������       �                     @        4       5                    :@�q�q�?             @        ������������������������       �                     �?        6       7                  S�2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        9       <                    �?z�G�z�?             $@       :       ;                 �&B@�<ݚ�?             "@       ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ?       `                    �?\�Uo��?             C@       @       Y                    �?<=�,S��?            �A@       A       N                    �?d��0u��?             >@       B       M                 ��&@p�ݯ��?             3@       C       J                 @3�@�t����?
             1@        D       G                 �?�@      �?              @        E       F                    9@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        H       I                   �8@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        K       L                    4@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        O       P                   �8@���|���?             &@        ������������������������       �                      @        Q       X                    C@�<ݚ�?             "@       R       W                   �@@�q�q�?             @       S       T                    ;@z�G�z�?             @        ������������������������       �                      @        U       V                 ��1@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        Z       _                 м�6@���Q��?             @       [       \                    <@�q�q�?             @        ������������������������       �                     �?        ]       ^                    @@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        a       b                    4@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        e       f                     @�\=lf�?+            �P@       ������������������������       �        *            �P@        ������������������������       �                     �?        ������������������������       �                     @        i       �                    �?���Ee�?6           p~@        j       �                  I>@R���Q�?1             T@       k       �                    �?�S����?#            �L@       l       �                 ��d5@�2����?"            �K@       m       �                 83�0@d}h���?             E@       n       q                   �6@:�&���?            �C@        o       p                 ��y@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        r       s                 ���@(N:!���?            �A@        ������������������������       �                     (@        t       w                     @�㙢�c�?             7@        u       v                 `��,@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        x                          �=@R���Q�?             4@       y       |                   @@z�G�z�?	             .@        z       {                   @<@����X�?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        }       ~                   �<@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �2@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     *@        ������������������������       �                      @        �       �                    �?�û��|�?             7@       �       �                    �?�d�����?             3@        �       �                 ��lK@����X�?             @        ������������������������       �                     �?        �       �                    �?r�q��?             @       ������������������������       �                     @        �       �                 �̾w@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                     �?      �?             (@       �       �                   �:@�z�G��?             $@        ������������������������       �                      @        �       �                   @H@      �?              @        �       �                 ���S@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    @�:�O�?           py@        �       �                    �?�q�q�?             5@        �       �                     @      �?              @       ������������������������       �                     @        �       �                    @      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                     @��
ц��?
             *@       ������������������������       �                     @        ������������������������       �                     @        �       .                  �R@åI$`�?�             x@       �       �                     �?     |�?�             x@        �       �                    �?�q�q�?/             R@        ������������������������       �                     �?        �       �                   �I@@���?T�?.            �Q@       �       �                    �?���!pc�?$            �K@       �       �                   �>@������?#             K@        �       �                   `G@D�n�3�?             3@       �       �                   �E@b�2�tk�?             2@       �       �                 ��$:@j���� �?             1@        ������������������������       �                     @        �       �                    @@�z�G��?             $@       �       �                   @>@և���X�?             @       �       �                 `fF<@      �?             @        ������������������������       �      �?             @        �       �                   �<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �;@b�h�d.�?            �A@        �       �                    7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 03�U@      �?             @@       �       �                    �? ��WV�?             :@       ������������������������       �        	             ,@        �       �                   �@@�8��8��?             (@        �       �                 `f�N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             0@        �       -                   �?4��?�?�            �s@       �                          �?L��B�?�            �q@       �                       0��D@�.�?�P�?�             n@       �       �                    �?�e)���?�            �m@        �       �                  ��@`2U0*��?             9@        ������������������������       �                     .@        �       �                 ��(@ףp=
�?	             $@       �       �                    >@      �?              @        �       �                   �<@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �                         �N@��-#���?�            �j@       �       �                 ���@Lő����?�            `j@        �       �                 �&b@�S����?             3@       �       �                 ���@�IєX�?             1@       ������������������������       �                     (@        �       �                 ��@z�G�z�?             @        �       �                    B@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   �?@�8��8N�?z             h@       �       �                     @P�2E��?S            @`@        �       �                    &@ 7���B�?             ;@        �       �                   �5@r�q��?             @        �       �                   �1@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     5@        �       �                 @3�@X�?٥�?A            �Y@        ������������������������       �                     �H@        �       �                   �<@h�WH��?!             K@       �       �                   �0@Hm_!'1�?            �H@        �       �                 pFD!@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 @3"@Du9iH��?            �E@       �       �                   �2@ �Cc}�?             <@        ������������������������       �                     @        �       �                 ��) @؇���X�?             5@       �       �                   �4@�X�<ݺ?             2@        ������������������������       �      �?              @        ������������������������       �        
             0@        �       �                    8@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        	             .@        �       �                 ���"@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?                               @3�@��� ��?'             O@                              �Y5@      �?             4@        ������������������������       �                      @              
                   E@�q�q�?
             (@                                A@�q�q�?             "@                                �@      �?             @        ������������������������       �                      @        ������������������������       �                      @              	                �?�@z�G�z�?             @       ������������������������       �                     @        ������������������������       �      �?              @                              P�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                @A@@4և���?             E@                                �@@@�0�!��?             1@        ������������������������       �                     @                              ��%@      �?             (@        ������������������������       �                     @        ������������������������       ����Q��?             @        ������������������������       �                     9@        ������������������������       �                     �?        ������������������������       �                     @                                   @&^�)b�?            �E@                                �7@      �?	             0@        ������������������������       �                     @                                 <@���|���?             &@        ������������������������       �                      @                                 �?X�<ݚ�?             "@                                C@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        !      $                   5@PN��T'�?             ;@        "      #                �Y�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        %      *                   �?�8��8��?             8@       &      )                  �9@      �?
             0@        '      (                  �8@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     *@        +      ,                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     =@        ������������������������       �                      @        �t�bh�h*h-K ��h/��R�(KM/KK��h]�B�        }@      o@      L@      e@      ,@      (@              @      ,@       @      @      @      @      @      �?               @      @              @       @      @               @       @      �?              �?       @              @               @      �?              �?       @              E@     �c@      B@     �c@     �A@     �V@     �A@     �U@              *@     �A@     @R@      @      D@      @      @      @      �?              �?      @                       @      �?     �B@              :@      �?      &@      �?       @      �?                       @              "@      ?@     �@@       @      2@      @      �?      �?      �?      �?                      �?       @              @      1@      @      ,@      @      @       @              �?      @              @      �?       @              �?      �?      �?      �?                      �?       @       @       @      @       @      @              @              �?              @      7@      .@      6@      *@      3@      &@      (@      @      (@      @      @      @      @      �?              �?      @              �?      @      �?                      @       @      �?              �?       @                       @      @      @               @      @       @      @       @      @      �?       @               @      �?              �?       @                      �?      @              @       @      �?       @              �?      �?      �?      �?                      �?       @              �?       @      �?                       @              @      �?     �P@             �P@      �?              @             �y@     �S@      O@      2@      H@      "@      G@      "@     �@@      "@      @@      @      �?      @      �?                      @      ?@      @      (@              3@      @       @      �?              �?       @              1@      @      (@      @      @       @      @       @      �?              @      �?      @                      �?      @              �?       @      �?                       @      *@               @              ,@      "@      ,@      @      @       @              �?      @      �?      @              �?      �?      �?                      �?      "@      @      @      @               @      @      �?       @      �?              �?       @              @               @                      @     �u@     �N@      @      ,@      �?      @              @      �?      @              @      �?              @      @              @      @             0u@     �G@     0u@     �F@     �L@      .@      �?              L@      .@      D@      .@      D@      ,@      &@       @      &@      @      $@      @      @              @      @      @      @      @      @       @       @      �?      �?              �?      �?                      �?              @      �?                      �?      =@      @      �?       @      �?                       @      <@      @      9@      �?      ,@              &@      �?      �?      �?              �?      �?              $@              @      @              @      @                      �?      0@             �q@      >@     �o@      >@     @k@      6@     @k@      3@      8@      �?      .@              "@      �?      @      �?       @      �?       @                      �?      @               @             @h@      2@     @h@      1@      0@      @      0@      �?      (@              @      �?      �?      �?              �?      �?              @                       @     @f@      ,@      _@      @      :@      �?      @      �?       @      �?      �?              �?      �?      @              5@             �X@      @     �H@             �H@      @     �F@      @      @      �?              �?      @              D@      @      9@      @      @              2@      @      1@      �?      �?      �?      0@              �?       @      �?                       @      .@              @      �?      @                      �?      K@       @      .@      @       @              @      @      @      @       @       @               @       @              @      �?      @              �?      �?      �?       @      �?                       @     �C@      @      ,@      @      @              "@      @      @               @      @      9@                      �?              @     �A@       @      (@      @      @              @      @       @              @      @       @      @              @       @              @              7@      @      �?       @      �?                       @      6@       @      .@      �?       @      �?       @                      �?      *@              @      �?              �?      @              =@                       @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ��DphG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMKhuh*h-K ��h/��R�(KMK��h|�B�R         �                    �?���x�W�?�           @�@               q                    @
��l۹�?�             o@              ^                   �>@D�4����?�            �k@                                   @�J��%�?c            `b@                                   �?���C��?%            �J@        ������������������������       �                     &@                                   �?؇���X�?             E@                                 �;@�t����?             A@       	                           �?z�G�z�?             4@       
                            �?�<ݚ�?             2@        ������������������������       �                     @                                   �?�q�q�?	             (@                                  �?X�<ݚ�?             "@                                  �6@      �?             @       ������������������������       �                     @        ������������������������       �                     @                                  �7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     ,@                                    �?      �?              @        ������������������������       �                      @        ������������������������       �                     @               9                    �?��V�I��?>            �W@               &                    �?����X�?             E@               !                    �?������?             .@                                    �?և���X�?             @                               ���%@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        "       %                    5@      �?              @        #       $                 83�0@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        '       8                    �?l��
I��?             ;@       (       )                    1@R�}e�.�?             :@        ������������������������       �                      @        *       7                    �?�q�q�?             8@       +       ,                    4@8����?             7@        ������������������������       �                     �?        -       .                 ���@���!pc�?             6@        ������������������������       �                      @        /       0                    9@z�G�z�?
             4@        ������������������������       �                      @        1       6                 pF @�<ݚ�?	             2@       2       3                 ���@      �?             0@        ������������������������       �                     @        4       5                 �&B@8�Z$���?             *@       ������������������������       �"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        :       A                    @
j*D>�?#             J@        ;       @                    �?؇���X�?             @       <       ?                    �?      �?             @       =       >                   �&@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        B       ]                    @�L�lRT�?            �F@       C       V                    �?���|���?             F@       D       U                    �?�q�q�?             >@       E       F                 ���@��}*_��?             ;@        ������������������������       �                     @        G       H                   �5@�q�q�?             8@        ������������������������       �                     @        I       J                   �@p�ݯ��?             3@        ������������������������       �                      @        K       P                 �]*@�t����?             1@       L       M                    :@�C��2(�?             &@        ������������������������       �                     @        N       O                   �;@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        Q       T                    ;@�q�q�?             @        R       S                    9@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        W       \                    �?և���X�?             ,@        X       Y                    �?؇���X�?             @        ������������������������       �                     @        Z       [                    1@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        _       h                 `f$@$G$n��?0            �R@        `       g                    �?�q�q�?             @       a       b                 ��n @      �?             @        ������������������������       �                     �?        c       d                  SE"@�q�q�?             @        ������������������������       �                     �?        e       f                    I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        i       j                     @l��\��?+             Q@       ������������������������       �        %            �M@        k       p                    C@�q�q�?             "@        l       o                   �@@      �?             @       m       n                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        r                           =@      �?             <@       s       t                    �?�<ݚ�?             ;@        ������������������������       �                     "@        u       ~                 ���d@�q�q�?             2@       v       }                   �6@z�G�z�?	             .@       w       x                    @�q�q�?             "@        ������������������������       �                     @        y       |                    @���Q��?             @       z       {                    @      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                 �?�@�.��q�?!           �|@        �       �                   @@@�\�)G�?Z            �`@       �       �                 �{@=�Ѝ;�?H            �Y@       �       �                    �?z���=��?7            @S@       �       �                    �?��A��?5            �R@       �       �                 ���@8�Z$���?0            @P@       �       �                    �?Du9iH��?            �E@        �       �                    5@ףp=
�?             4@        �       �                 �{@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ���@�X�<ݺ?             2@        ������������������������       �                     @        �       �                   @<@�8��8��?             (@       �       �                    9@r�q��?             @        ������������������������       �                     �?        ������������������������       �z�G�z�?             @        ������������������������       �                     @        �       �                    7@�nkK�?             7@        ������������������������       �                     &@        �       �                 �&b@�8��8��?
             (@       ������������������������       �                     @        �       �                 ���@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 P�N@�X����?             6@       �       �                 �1@�E��ӭ�?             2@       �       �                   �3@�t����?             1@        ������������������������       �                      @        �       �                 ��@�q�q�?             .@        �       �                   �>@      �?              @       �       �                   �<@�q�q�?             @       ������������������������       �z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 �?$@և���X�?             @        ������������������������       �      �?              @        �       �                   �;@���Q��?             @       �       �                   �6@�q�q�?             @        ������������������������       �                     �?        �       �                   �9@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                    :@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �7@�q�q�?             "@        ������������������������       �                     @        �       �                   �9@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     :@        ������������������������       �                     @@        �       �                     �?�A����?�            �t@        �       �                    �?�qs�_�?:            �Z@       �       �                    @��H���?8            @Y@       �       �                   �1@�fSO��?7            �X@        ������������������������       �                     @        �       �                   �8@$)}�~z�?5            �W@        ������������������������       �                     @        �       �                    �? 9�����?1             V@       �       �                   �?@��
ц��?%            @P@       �       �                 `f�B@p�ݯ��?             C@       �       �                   �<@
;&����?             7@       �       �                    �?ҳ�wY;�?
             1@        �       �                 �ܵ<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 `fF:@X�Cc�?             ,@        ������������������������       �                      @        �       �                   �;@      �?             (@        ������������������������       �                      @        �       �                 `fF<@�z�G��?             $@        ������������������������       ����Q��?             @        �       �                   �>@z�G�z�?             @        ������������������������       �                     @        �       �                   �@@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?z�G�z�?	             .@        �       �                   �;@      �?              @        �       �                    �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                   @B@�5��?             ;@        �       �                   �A@�8��8��?             (@        ������������������������       �                     @        �       �                 @�Cq@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �?@�q�q�?             .@       �       �                    �?����X�?             @        ������������������������       �                     �?        �       �                   @G@r�q��?             @        �       �                 03k:@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?
;&����?             7@       �       �                    ;@և���X�?             5@        ������������������������       �                     @        �       �                   �F@�q�q�?
             2@        ������������������������       �                      @        �       �                 @�pX@���Q��?             $@       �       �                   @P@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       8                   �?�����?�            �k@       �       1                   �?n�3���?b             c@       �       0                  �F@��f/w�?M            �^@       �       )                  �B@�n����?C            @Z@       �                          �?�n`���?=            @W@        �       �                 �R,@      �?              @        ������������������������       �                      @        �       �                     @r�q��?             @        ������������������������       �                     �?                               `v�0@z�G�z�?             @        ������������������������       �                      @                                �2@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                  @@�0�!��?8            @U@              	                  �5@@�0�!��?             1@                                 &@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        
                        �'@�8��8��?	             (@        ������������������������       �                     @                                �>@؇���X�?             @       ������������������������       �                     @        ������������������������       �      �?              @                                �0@@�0�!��?+             Q@        ������������������������       ��q�q�?             @              (                  @@@8�Z$���?)            @P@                             ��i @"pc�
�?$            �K@                               �3@r֛w���?             ?@        ������������������������       ����Q��?             @                                 ;@���B���?             :@        ������������������������       �                     @                                 ?@      �?             4@                                =@������?
             1@                             ��) @      �?	             0@       ������������������������       �                     (@        ������������������������       �                     @        ������������������������       �                     �?                              @3�@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?               %                  �<@�8��8��?             8@       !      "                �T�C@���7�?             6@       ������������������������       �                     2@        #      $                   ;@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        &      '                ���"@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        *      -                    @�q�q�?             (@        +      ,                  @D@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        .      /                ��	0@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             1@        2      3                    @(;L]n�?             >@        ������������������������       �                     (@        4      7                   �?�X�<ݺ?             2@       5      6                  �6@�8��8��?
             (@        ������������������������       �                     �?        ������������������������       �        	             &@        ������������������������       �                     @        9      D                   �?ٜSu��?+            @Q@       :      C                   @���|���?             F@       ;      >                03{3@�g�y��?             ?@        <      =                   ?@$�q-�?             *@       ������������������������       �                     (@        ������������������������       �                     �?        ?      @                039@�<ݚ�?             2@        ������������������������       �                      @        A      B                   +@���Q��?	             $@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     *@        E      F                   �?H%u��?             9@        ������������������������       �                     �?        G      J                   @�8��8��?             8@        H      I                   @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     5@        �t�bh�h*h-K ��h/��R�(KMKKK��h]�B�       P{@     0q@     �S@     @e@      M@     `d@      H@     �X@      @     �G@              &@      @      B@      @      >@      @      0@      @      ,@              @      @       @      @      @      @      @              @      @              �?       @      �?                       @              @               @              ,@       @      @       @                      @      E@      J@      (@      >@      @      &@      @      @       @      @              @       @              �?              �?      @      �?      @      �?                      @              @       @      3@      @      3@               @      @      1@      @      0@      �?              @      0@       @              @      0@               @      @      ,@       @      ,@              @       @      &@       @      "@               @       @                      �?      �?              >@      6@      �?      @      �?      @      �?       @      �?                       @              �?              @      =@      0@      <@      0@      4@      $@      1@      $@              @      1@      @      @              (@      @               @      (@      @      $@      �?      @              @      �?              �?      @               @      @       @      �?              �?       @                      @      @               @      @      �?      @              @      �?       @      �?                       @      @              �?              $@      P@      @       @       @       @      �?              �?       @              �?      �?      �?      �?                      �?       @              @      O@             �M@      @      @      �?      @      �?       @      �?                       @              �?      @              5@      @      5@      @      "@              (@      @      (@      @      @      @      @               @      @      �?      @      �?                      @      �?              @                      @              �?     `v@     @Z@     �^@      *@     �V@      *@      P@      *@     �N@      *@     �K@      $@      D@      @      2@       @      �?      �?      �?                      �?      1@      �?      @              &@      �?      @      �?      �?              @      �?      @              6@      �?      &@              &@      �?      @              @      �?              �?      @              .@      @      *@      @      (@      @       @              $@      @      @       @      @       @      @      �?              �?       @              @      @      �?      �?      @       @      �?       @              �?      �?      �?      �?                      �?       @              �?               @       @       @                       @      @      @      @               @      @              @       @              @              :@              @@             �m@      W@     �N@      G@     �K@      G@     �J@      G@              @     �J@     �D@      @             �G@     �D@     �A@      >@      8@      ,@      (@      &@      @      &@      �?       @      �?                       @      @      "@       @              @      "@               @      @      @       @      @      �?      @              @      �?      �?      �?                      �?      @              (@      @      @      @       @      @              @       @              @              @              &@      0@      �?      &@              @      �?      @      �?                      @      $@      @       @      @      �?              �?      @      �?      �?              �?      �?                      @       @              (@      &@      (@      "@              @      (@      @       @              @      @      �?      @              @      �?              @                       @       @              @             �e@      G@     @_@      ;@      X@      :@     �S@      :@     �R@      2@      @      @               @      @      �?      �?              @      �?       @               @      �?       @                      �?     �Q@      .@      ,@      @      @       @               @      @              &@      �?      @              @      �?      @              �?      �?      L@      (@      �?       @     �K@      $@     �F@      $@      7@       @       @      @      5@      @      @              .@      @      *@      @      (@      @      (@                      @      �?               @      �?       @                      �?      6@       @      5@      �?      2@              @      �?              �?      @              �?      �?      �?                      �?      $@              @       @      @      �?      �?               @      �?      �?      @              @      �?              1@              =@      �?      (@              1@      �?      &@      �?              �?      &@              @              I@      3@      <@      0@      .@      0@      �?      (@              (@      �?              ,@      @       @              @      @              @      @              *@              6@      @              �?      6@       @      �?       @               @      �?              5@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ%�[6hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B�G         L                    �?�25����?�           @�@                                    @�<ݚ�?�            @m@                                 �;@`���i��?P            �`@                                   �?t��ճC�?             F@        ������������������������       �        
             .@               	                     �?ܷ��?��?             =@                                   �?����X�?             @       ������������������������       �                     @        ������������������������       �                      @        
                          �9@���7�?             6@       ������������������������       �                     4@                                  �/@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        3             V@               %                    �?4�M�f��?F            �Y@               $                    @      �?             B@              !                    �?�������?             A@                                  �?V�a�� �?             =@                                 �+@�J�4�?             9@                                  2@      �?             8@        ������������������������       �                     @                                   �?r�q��?             2@        ������������������������       �                     �?                                  �5@@�0�!��?             1@        ������������������������       �                     �?                                ���@      �?
             0@        ������������������������       �                      @        ������������������������       �        	             ,@        ������������������������       �                     �?                                 ���.@      �?             @        ������������������������       �                      @        ������������������������       �                      @        "       #                    �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        &       '                 ���@����e��?-            �P@        ������������������������       �                     @        (       G                     @�e�,��?)            �M@       )       6                 `f�%@Z�K�D��?!            �G@       *       +                 �?�@�J�4�?             9@        ������������������������       �                     &@        ,       3                    �?����X�?             ,@       -       0                 @3�@      �?
             (@        .       /                   �8@      �?             @        ������������������������       �                      @        ������������������������       �                      @        1       2                   �I@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        4       5                   �#@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        7       D                    �?8�A�0��?             6@       8       C                   �@@z�G�z�?             .@       9       B                 `fV6@      �?	             (@       :       ;                 @3�,@"pc�
�?             &@        ������������������������       �                     @        <       =                    ;@      �?              @        ������������������������       �                     �?        >       ?                 ��1@؇���X�?             @        ������������������������       �                     @        @       A                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        E       F                    0@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        H       K                    @r�q��?             (@       I       J                    ,@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        M       x                 �?�@�NG�#=�?/           �}@        N       w                    �?,I�e���?\            �b@       O       p                 �1@��[�?Z            �b@       P       o                    =@8�Z$���?=             Z@       Q       R                   �3@6��f�?+            @S@        ������������������������       �                     @        S       V                   �5@\�CX�?&            �Q@        T       U                 P�@      �?              @        ������������������������       �                     @        ������������������������       �                     @        W       d                  ��@Z���c��?"            �O@       X       [                    �?�*/�8V�?            �G@        Y       Z                 ���@z�G�z�?             .@        ������������������������       �                     @        ������������������������       �      �?             (@        \       c                 ���@      �?             @@       ]       ^                   �8@�����H�?
             2@        ������������������������       �                     �?        _       b                   �;@�IєX�?	             1@        `       a                 ��@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        ������������������������       �                     ,@        e       h                    �?      �?
             0@        f       g                    �?      �?              @       ������������������������       �և���X�?             @        ������������������������       �                     �?        i       j                   �7@      �?              @        ������������������������       �                     �?        k       n                 �?$@����X�?             @       l       m                    �?���Q��?             @       ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     ;@        q       v                    �?`���i��?             F@        r       u                    @@      �?             @       s       t                   �<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     D@        ������������������������       �                     @        y       �                    �?�]N���?�            pt@        z       �                    �?�eP*L��?$            �K@       {       |                    @f���M�?             ?@        ������������������������       �                     @        }       ~                 �R,@����X�?             <@        ������������������������       �                      @               �                   �J@�θ�?             :@       �       �                 �̾w@�㙢�c�?             7@       �       �                    =@��2(&�?             6@       �       �                    �?     ��?             0@       �       �                     �?�θ�?	             *@       �       �                    9@      �?              @        ������������������������       �                     �?        �       �                 �ܵ<@����X�?             @        ������������������������       �                     @        �       �                 03SA@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �8@z�G�z�?             @        ������������������������       �                      @        �       �                    ;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                 ��L@@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�q�q�?             8@       �       �                 �U�X@�û��|�?             7@       �       �                   �9@�q�q�?             5@        ������������������������       �                     &@        �       �                    �?�z�G��?	             $@       �       �                 @3�J@      �?              @       ������������������������       �                     @        �       �                    C@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                     �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                    @l�]�NG�?�             q@        �       �                    �?�X����?             6@        ������������������������       �                     �?        �       �                    @����X�?             5@       ������������������������       �        	             *@        �       �                 ���A@      �?              @        �       �                 @3;:@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �                          @z�G�z�?�            @o@       �       �                 @3�@��[�p�?�            `m@        �       �                    �?��.k���?
             1@       �       �                   �D@�	j*D�?             *@       �       �                    �?���Q��?             $@       �       �                    :@X�<ݚ�?             "@        ������������������������       �                     �?        �       �                   �A@      �?              @       �       �                   �?@z�G�z�?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                     �?�	{���?�            @k@        �       �                    >@L
�q��?$            �M@        �       �                   �<@"pc�
�?             6@       �       �                   �;@����X�?             ,@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �>@      �?	             (@        �       �                 `fF<@���Q��?             @        ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                   �J@��J�fj�?            �B@       �       �                    �?X�<ݚ�?             ;@       �       �                 �T!@@���Q��?             9@        �       �                   �G@8�Z$���?             *@        �       �                    G@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �D@�q�q�?             (@        ������������������������       �                      @        �       �                   @H@z�G�z�?             $@       ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �?@ףp=
�?             $@       �       �                 `fF<@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    )@^�!~X�?k            �c@        ������������������������       �                     �?        �                          M@�+ت�M�?j            �c@       �                          �?�䞠�l�?h            @c@       �       �                   �0@��E�B��?`            �a@        �       �                 �̌"@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �                           @ ���g=�?^            @a@        �       �                    �?R���Q�?%             N@       �       �                   �*@�*/�8V�?            �G@       �       �                    ;@$G$n��?            �B@        ������������������������       �        	             .@        �       �                 `fF)@�GN�z�?             6@        ������������������������       �                     @        �       �                    =@�d�����?             3@        ������������������������       �                      @        �       �                    G@@�0�!��?
             1@       �       �                    @@      �?             (@        ������������������������       �                     @        �       �                   @D@      �?              @       �       �                   @B@�q�q�?             @       ������������������������       ����Q��?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     $@        �                          �@@�	j*D�?             *@        �       �                   �>@      �?              @        ������������������������       �                     @        �       �                   �H@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @                                @@@�:�^���?9            �S@                                �?�^����?-            �M@                                ?@ܷ��?��?,             M@                                �?�X�<ݺ?)             K@        ������������������������       �                     @                                 �?��<D�m�?%            �H@                             �T�C@@4և���?              E@       	                        �;@�}�+r��?             C@       
                        �:@�����?             5@                             ��Y @P���Q�?             4@                                 4@؇���X�?             @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �        	             *@        ������������������������       �                     �?        ������������������������       �                     1@        ������������������������       �      �?             @        ������������������������       �                     @                              ��i @      �?             @        ������������������������       �                      @                              d�6@@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     3@        ������������������������       �                     *@                                �P@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     .@        �t�b��;     h�h*h-K ��h/��R�(KMKK��h]�B�       pz@     r@      J@     �f@      @      `@      @     �D@              .@      @      :@       @      @              @       @              �?      5@              4@      �?      �?              �?      �?                      V@     �H@     �J@      "@      ;@      "@      9@      @      7@      @      5@      @      5@              @      @      .@              �?      @      ,@      �?               @      ,@       @                      ,@      �?               @       @       @                       @      @       @      @                       @               @      D@      :@              @      D@      3@      >@      1@      5@      @      &@              $@      @      "@      @       @       @       @                       @      @      �?      @                      �?      �?      �?              �?      �?              "@      *@      @      (@      @      "@       @      "@              @       @      @      �?              �?      @              @      �?       @      �?                       @      �?                      @      @      �?              �?      @              $@       @      @       @      @                       @      @             0w@     �Z@     �`@      1@     ``@      1@      V@      0@     �N@      0@      @             �K@      0@      @      @      @                      @      I@      *@      E@      @      (@      @      @              "@      @      >@       @      0@       @              �?      0@      �?      @      �?              �?      @              (@              ,@               @       @      @      @      @      @      �?              @      @      �?               @      @       @      @       @       @              �?               @      ;@             �E@      �?      @      �?      �?      �?      �?                      �?       @              D@              @             �m@     �V@      >@      9@      4@      &@              @      4@       @               @      4@      @      3@      @      3@      @      *@      @      $@      @      @       @      �?              @       @      @              �?       @               @      �?              @      �?       @               @      �?              �?       @              @              @                      �?      �?       @      �?                       @      $@      ,@      "@      ,@      @      ,@              &@      @      @      @       @      @              �?       @      �?                       @      �?      �?              �?      �?               @              �?             �i@     @P@      @      .@      �?              @      .@              *@      @       @       @       @       @                       @      @              i@      I@      g@      I@       @      "@      @      "@      @      @      @      @      �?              @      @      �?      @               @      �?       @       @      �?              �?              @      @              f@     �D@     �C@      4@      2@      @      $@      @      �?      �?              �?      �?              "@      @       @      @       @      �?               @      @               @              5@      0@      (@      .@      $@      .@       @      &@       @      @              @       @                       @       @      @               @       @       @      @               @       @       @                       @       @              "@      �?      @      �?      @                      �?      @             @a@      5@              �?     @a@      4@      a@      2@     �^@      2@      �?       @               @      �?             �^@      0@     �I@      "@      E@      @      @@      @      .@              1@      @      @              ,@      @               @      ,@      @      "@      @      @              @      @      @       @      @       @      �?              �?      �?      @              $@              "@      @      @      @      @              �?      @              @      �?              @             �Q@      @      J@      @      J@      @     �I@      @      @              G@      @     �C@      @      B@       @      3@       @      3@      �?      @      �?      �?      �?      @              *@                      �?      1@              @      �?      @              �?      @               @      �?      �?      �?                      �?              �?      3@              *@               @       @               @       @              .@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�	3 hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMChuh*h-K ��h/��R�(KMC��h|�B�P         �                 `f�%@T�����?�           @�@                                    �?.�*���?�            �r@        ������������������������       �                     @               	                 ���@�V���1�?�            �r@                                  �;@������?             B@                                   :@�IєX�?	             1@       ������������������������       �                     0@        ������������������������       �                     �?        ������������������������       �        
             3@        
       #                   �4@ά��.��?�            @p@                                   �?*O���?             B@                                ���@z�G�z�?             @        ������������������������       �                     @                                   ,@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               "                    �?¦	^_�?             ?@                                  �?������?             >@                                  �?���B���?             :@                                03�@�q�q�?             @        ������������������������       �                     �?                                   0@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?                                   1@R���Q�?             4@                                �̌!@�<ݚ�?             "@        ������������������������       ��q�q�?             @        ������������������������       �                     @                                    @�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@                !                    3@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        $       �                    �?d}h���?�             l@       %       &                 ��@0ݪ��?�            �k@        ������������������������       �                     �?        '       �                   @N@��t��\�?�            �k@       (       }                 @3�@�{��?��?�             k@       )       t                   @@@,A����?\            �b@       *       k                   �>@�&�5y�?N             _@       +       ^                 �̌@4և����?G             \@       ,       =                    �?����X�?2            @S@        -       .                   �5@�<ݚ�?             2@        ������������������������       �                     �?        /       0                    �?@�0�!��?             1@        ������������������������       �                     �?        1       2                    8@     ��?             0@        ������������������������       �                     @        3       4                   �9@�θ�?
             *@        ������������������������       �                     �?        5       <                    �?r�q��?	             (@       6       ;                    �?�C��2(�?             &@       7       :                 �&B@ףp=
�?             $@       8       9                 ���@؇���X�?             @        ������������������������       �                      @        ������������������������       �z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        >       W                    �?(2��R�?$            �M@       ?       H                    �?0��_��?             �J@        @       C                 ���@r�q��?	             (@        A       B                   �7@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        D       E                    9@      �?              @        ������������������������       �                      @        F       G                   @<@r�q��?             @       ������������������������       �z�G�z�?             @        ������������������������       �                     �?        I       N                   �5@��p\�?            �D@        J       K                 @�@����X�?             @        ������������������������       �                     @        L       M                 ��L@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        O       P                    �?г�wY;�?             A@        ������������������������       �                     .@        Q       R                 �?$@�}�+r��?             3@       ������������������������       �                     .@        S       T                   �9@      �?             @        ������������������������       �                      @        U       V                   �;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        X       Y                    �?      �?             @        ������������������������       �                     �?        Z       [                   �7@���Q��?             @        ������������������������       �                     �?        \       ]                   �9@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        _       d                 �?�@(N:!���?            �A@       `       c                    �? ��WV�?             :@        a       b                   �<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     8@        e       j                    �?�q�q�?             "@       f       i                    �?և���X�?             @       g       h                    9@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        l       m                 �&B@�q�q�?             (@        ������������������������       �                      @        n       o                   �?@z�G�z�?             $@        ������������������������       �                     @        p       q                   �@����X�?             @        ������������������������       �                      @        r       s                 �?�@���Q��?             @        ������������������������       �                     �?        ������������������������       �      �?             @        u       v                    �?ȵHPS!�?             :@        ������������������������       �                     @        w       x                    �?؇���X�?
             5@        ������������������������       �                     @        y       z                 �?�@     ��?	             0@       ������������������������       �                     (@        {       |                   �D@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ~                        `�X!@��IF�E�?.            �P@        ������������������������       �                    �A@        �       �                 ��!@��a�n`�?             ?@        ������������������������       �                      @        �       �                     @д>��C�?             =@        �       �                    �?�q�q�?	             (@        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�IєX�?             1@        ������������������������       �                     $@        �       �                   �<@؇���X�?             @       ������������������������       �                     @        �       �                   �"@�q�q�?             @        ������������������������       �                     �?        �       �                    ?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ��\!@      �?             @        ������������������������       �                      @        �       �                     @      �?             @       �       �                   �P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?\����?�            �y@        �       �                    @�j��e�?u            �f@       �       �                     @pc�
��?q             f@       �       �                   �;@$Q�q�?M            �_@        �       �                    6@؇���X�?             E@        �       �                   �1@X�<ݚ�?             "@       �       �                 ��*@�q�q�?             @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                 ���`@Pa�	�?            �@@       ������������������������       �                     >@        �       �                 03�g@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �H@�Ń��̧?1             U@       ������������������������       �        (            �Q@        �       �                   @I@؇���X�?	             ,@        �       �                 03[;@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     $@        �       �                    �?z�):���?$             I@        �       �                 ��.@ҳ�wY;�?             1@        �       �                    �?      �?              @       �       �                    �?����X�?             @        ������������������������       �                     @        �       �                 P��+@      �?             @        ������������������������       �                     �?        �       �                    �?�q�q�?             @        ������������������������       �                     �?        �       �                   �<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        �       �                     @�'�=z��?            �@@       �       �                   �D@�X����?             6@       �       �                    �?      �?             4@        �       �                    1@�����H�?             "@        �       �                 `f7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �@@���|���?	             &@       �       �                 ���5@X�<ݚ�?             "@       �       �                    �?      �?              @        �       �                   �=@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 P��)@      �?             @        ������������������������       �                     �?        �       �                   �=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                   �>@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                     @        �       B                  �R@�D�>��?�            �l@       �       7                Ј�V@     ��?�             l@       �                          �?�E���?            �i@       �                          �?2%ޑ��?Y            �a@       �                           @���>���?V            �`@       �       �                    :@pN�Z��?C            �Z@        ������������������������       �                     ;@        �       �                     �?     ��?6             T@       �       �                 Ј�U@��[�8��?!            �I@       �       �                   �>@z�G�z�?              I@        �       �                    ?@�X����?             6@        �       �                 ���<@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        �       �                    �?      �?	             (@        �       �                   �F@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ��:@X�<ݚ�?             "@        ������������������������       �                     �?        �       �                 `f�<@      �?              @       �       �                   �K@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                   �J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 8�<Q@ �Cc}�?             <@       �       �                    @@���N8�?             5@       �       �                 `f�B@ףp=
�?             $@        �       �                   �A@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        �       �                    �?����X�?             @        ������������������������       �                     �?        �       �                   @G@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?                                 �E@\-��p�?             =@                               @C@      �?             0@                                �?؇���X�?             ,@                                �?ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@                                 �?      �?             @        ������������������������       �                     �?              	                  �>@�q�q�?             @        ������������������������       �                     �?        
                        �@@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     *@                                 �?R�}e�.�?             :@                                 3@      �?             @        ������������������������       �                     �?                                 �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                 �?"pc�
�?             6@                             �T)D@������?	             .@       ������������������������       �                      @                                 ;@և���X�?             @        ������������������������       �                     �?                                 >@      �?             @       ������������������������       ����Q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @              &                   �?��&����?&            @P@               !                ���6@�eP*L��?             &@        ������������������������       �                     @        "      #                   �?r�q��?             @        ������������������������       �                     @        $      %                   �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        '      2                   �?�{��?��?!             K@       (      )                   �?����>�?            �B@        ������������������������       �                     @        *      -                   :@�4�����?             ?@        +      ,                   $@     ��?
             0@       ������������������������       �                     "@        ������������������������       �                     @        .      1                   &@��S�ۿ?
             .@        /      0                  C@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        3      6                   @�IєX�?             1@        4      5                   +@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        8      A                   @�\��N��?
             3@       9      @                  �L@      �?	             0@       :      ?                `f�e@����X�?             ,@       ;      >                �y[@�C��2(�?             &@        <      =                �U�X@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �t�bh�h*h-K ��h/��R�(KMCKK��h]�B0       0|@     Pp@      n@      O@      @             @m@      O@     �A@      �?      0@      �?      0@                      �?      3@             �h@     �N@      7@      *@      �?      @              @      �?      �?              �?      �?              6@      "@      6@       @      5@      @      @       @              �?      @      �?      @                      �?      1@      @      @       @      �?       @      @              $@      �?              �?      $@              �?      @      �?                      @              �?      f@      H@     �e@      H@              �?     �e@     �G@     �e@      F@     @\@     �B@     �V@      A@     �U@      :@     �K@      6@      @      ,@      �?              @      ,@              �?      @      *@              @      @      $@      �?               @      $@      �?      $@      �?      "@      �?      @               @      �?      @              @              �?      �?             �I@       @      H@      @      $@       @      @      �?              �?      @              @      �?       @              @      �?      @      �?      �?              C@      @      @       @      @              �?       @               @      �?             �@@      �?      .@              2@      �?      .@              @      �?       @              �?      �?              �?      �?              @      @      �?               @      @      �?              �?      @              @      �?              ?@      @      9@      �?      �?      �?      �?                      �?      8@              @      @      @      @      @      @      @                      @      �?               @              @       @       @               @       @              @       @      @               @       @      @      �?              �?      @      7@      @      @              2@      @      @              *@      @      (@              �?      @      �?                      @     �M@      @     �A@              8@      @               @      8@      @       @      @              @       @              0@      �?      $@              @      �?      @               @      �?      �?              �?      �?              �?      �?              @      @       @              �?      @      �?      �?              �?      �?                       @      �?             `j@     �h@      B@      b@      ?@      b@       @     �]@      @      B@      @      @       @      @       @      �?              �?       @                      @      @              �?      @@              >@      �?       @      �?                       @       @     �T@             �Q@       @      (@       @       @               @       @                      $@      7@      ;@      @      &@      @       @      @       @      @               @       @              �?       @      �?      �?              �?      �?      �?                      �?      �?                      "@      1@      0@      @      .@      @      .@      �?       @      �?       @               @      �?                      @      @      @      @      @      @      @      �?      @              @      �?               @       @              �?       @      �?       @                      �?      �?                       @       @              $@      �?      $@                      �?      @             �e@      K@     �e@     �H@     �d@     �C@     �]@      6@     �[@      6@      W@      .@      ;@             @P@      .@      D@      &@      D@      $@      .@      @      "@      �?      "@                      �?      @      @       @      �?              �?       @              @      @      �?              @      @       @      @              @       @              �?      �?              �?      �?              9@      @      4@      �?      "@      �?      @      �?      @                      �?      @              &@              @       @              �?      @      �?      @                      �?              �?      9@      @      (@      @      (@       @      "@      �?              �?      "@              @      �?      �?               @      �?      �?              �?      �?              �?      �?                       @      *@              3@      @      �?      @              �?      �?       @               @      �?              2@      @      &@      @       @              @      @              �?      @      @      @       @              �?      @              @              H@      1@      @      @              @      @      �?      @               @      �?              �?       @             �E@      &@      ;@      $@      @              5@      $@      @      "@              "@      @              ,@      �?      @      �?              �?      @              $@              0@      �?      @      �?              �?      @              "@              "@      $@      @      $@      @      $@      �?      $@      �?      @              @      �?                      @      @               @              @                      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ��.hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMmhuh*h-K ��h/��R�(KMm��h|�B@[                             @(����7�?�           @�@               	                     @�q�q�?            �C@                                   �?�����H�?             ;@                                   �?և���X�?             @        ������������������������       �                      @                                   �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     4@        
                           @r�q��?             (@       ������������������������       �                     @                                   �?���Q��?             @        ������������������������       �                      @                                ��T?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @               �                   �<@���v��?�           �@              =                     �?�~�#�?
           �z@               ,                    �?^��>�b�?'            @P@              %                    �?�`���?            �H@                               ��M@�Q����?             D@                                  �?�X����?             6@        ������������������������       �                     @                                  �>@j���� �?
             1@                                  �?�z�G��?             $@        ������������������������       �                      @                                   <@      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @                                    �?�<ݚ�?             2@       ������������������������       �                     &@        !       $                   �;@և���X�?             @       "       #                 ���Z@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        &       '                    3@X�<ݚ�?             "@        ������������������������       �                     @        (       )                    �?r�q��?             @        ������������������������       �                      @        *       +                   �8@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        -       8                 03�a@      �?             0@       .       7                    �?8�Z$���?
             *@       /       2                 0�"K@z�G�z�?	             $@        0       1                    7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        3       4                    �?      �?              @       ������������������������       �                     @        5       6                 �U�X@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        9       <                    �?�q�q�?             @       :       ;                   �5@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        >       �                    @\O�΄��?�            �v@       ?       �                 �%@��Q���?�            �v@       @       O                   �2@�^���?�             k@        A       D                    /@     ��?             @@        B       C                    �?�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        E       F                    �?$��m��?             :@        ������������������������       �                     �?        G       H                    �?`�Q��?             9@        ������������������������       �                     @        I       N                   �0@�KM�]�?	             3@        J       M                 �̌"@      �?              @       K       L                 pf�@���Q��?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     &@        P       �                 ���@��G���?v             g@       Q       R                   �4@�����?A            �W@        ������������������������       �                     "@        S       h                    �?8�$�>�?;            �U@        T       U                 �&�@������?             ;@        ������������������������       �                     @        V       g                    �?�q�q�?             8@       W       b                    �?�GN�z�?             6@       X       Y                   �5@�<ݚ�?             2@        ������������������������       �                     �?        Z       [                  ��@@�0�!��?
             1@        ������������������������       �                      @        \       ]                    9@��S�ۿ?	             .@        ������������������������       �                     �?        ^       a                 �&B@@4և���?             ,@       _       `                 ���@�8��8��?             (@        ������������������������       �                     �?        ������������������������       ��C��2(�?             &@        ������������������������       �                      @        c       d                 ���@      �?             @        ������������������������       �                      @        e       f                   �9@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        i       �                    �?�:�B��?)            �M@       j       {                    �?�2����?%            �K@       k       p                   �7@��� ��?             ?@        l       m                   �5@      �?              @        ������������������������       �                      @        n       o                 ���@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        q       r                 ���@���}<S�?             7@        ������������������������       �                     @        s       v                    �?�KM�]�?             3@        t       u                   @<@r�q��?             @       ������������������������       �z�G�z�?             @        ������������������������       �                     �?        w       x                  ��@$�q-�?	             *@        ������������������������       �                     @        y       z                 ��(@�����H�?             "@       ������������������������       �r�q��?             @        ������������������������       �                     @        |       }                     @�q�q�?             8@        ������������������������       �                     @        ~       �                   �5@      �?             4@               �                  s@      �?             @        ������������������������       �                     �?        �       �                 �1@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �:@     ��?             0@       �       �                 ���@�8��8��?             (@        �       �                   �8@z�G�z�?             @        �       �                 ���@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   �;@      �?             @        ������������������������       �                     �?        �       �                 pf�@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                 ��@      �?             @        ������������������������       �                      @        �       �                   �9@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                     @�X�<ݺ?5            �V@        �       �                    �?      �?              @        ������������������������       �                     �?        �       �                   �5@؇���X�?             @        ������������������������       ��q�q�?             @        ������������������������       �                     @        �       �                    �?Ћ����?0            �T@        �       �                    �?�����H�?             "@       �       �                 @3�@؇���X�?             @        �       �                   �8@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?��pBI�?)            @R@        ������������������������       �                     �?        �       �                   �4@������?(             R@        �       �                    �?�<ݚ�?             "@       �       �                   �3@      �?              @       �       �                 `�8"@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        "            �O@        �       �                    @x�f��^�?Y            �a@       �       �                   �7@��Zy�?J            @]@        �       �                 �&@�^�����?            �E@        ������������������������       �                     @        �       �                    �?�θ�?            �C@       �       �                    �?�J�4�?             9@       �       �                   �4@�}�+r��?             3@       ������������������������       �                     &@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                      @        �       �                 0339@      �?             @        �       �                 03�7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?X�Cc�?
             ,@        ������������������������       �                     @        �       �                 03�0@"pc�
�?             &@        �       �                    .@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�����H�?             "@       �       �                   �2@z�G�z�?             @        ������������������������       �                     @        �       �                   0>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �8@��+��?.            �R@        �       �                    �?8�Z$���?             *@       �       �                   �+@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        �       �                     @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �=@�p����?'            �N@       �       �                   �;@���Q��?#            �K@        �       �                    �?�㙢�c�?             7@        ������������������������       �                     @        �       �                   �9@P���Q�?             4@       �       �                    �?�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     &@        �       �                 `ff+@     ��?             @@        ������������������������       �                      @        �       �                    �?�q�q�?             8@        �       �                    �?"pc�
�?             &@        ������������������������       �                      @        �       �                 pF�-@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?$�q-�?             *@       �       �                    �?      �?              @       ������������������������       �                     @        �       �                  �v6@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    ;@r�q��?             @        ������������������������       �                      @        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     :@        ������������������������       �                     @        �       F                    @V�s�s�?�            �n@       �       =                03?U@�o;����?l            �c@       �       $                  @I@      �?[            �`@       �       #                 �}S@(옄��??             W@       �                         �G@~�4_�g�?=             V@       �                          �?`��_��?4            �Q@       �       �                    �?�>$�*��?            �D@        ������������������������       �                     *@        �                           �?�>4և��?             <@        �       �                   @E@r�q��?             (@       ������������������������       �                     @                               `f?@����X�?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?                                �@@     ��?             0@        ������������������������       �                     @                                 �?���!pc�?	             &@                                ,@�z�G��?             $@             
                  @D@և���X�?             @             	                  @A@�q�q�?             @       ������������������������       �      �?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?                                 �?���Q��?             >@        ������������������������       �                     *@                                 �?�t����?             1@                               �@@     ��?             0@                                 �?և���X�?             @        ������������������������       �                     �?                                 :@�q�q�?             @        ������������������������       �                      @                                @K@      �?             @       ������������������������       �                      @        ������������������������       �                      @                                  �?�����H�?             "@                                 �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?                                  �?@�0�!��?	             1@       ������������������������       �                     "@        !      "                  �H@      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        %      &                   �?�D����?             E@        ������������������������       �        	             (@        '      8                    �?r�q��?             >@       (      3                   �?�<ݚ�?             2@       )      2                   @@z�G�z�?	             .@       *      -                `fF<@      �?              @        +      ,                  @L@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        .      /                  @>@      �?             @        ������������������������       �                     �?        0      1                  �J@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        4      5                   L@�q�q�?             @        ������������������������       �                     �?        6      7                  @P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        9      <                   �?�8��8��?             (@       :      ;                  @N@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        >      ?                   �?      �?             8@       ������������������������       �        
             .@        @      E                   �?�q�q�?             "@       A      B                @�pX@և���X�?             @        ������������������������       �                      @        C      D                @�ys@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        G      L                   �?RB)��.�?6            �U@        H      I                   �?�eP*L��?             &@        ������������������������       �                     �?        J      K                   ?@���Q��?             $@        ������������������������       �                     @        ������������������������       �                     @        M      l                   @�7�QJW�?1            �R@       N      O                   �?�����?-             Q@        ������������������������       �                     @        P      e                   �?     ��?*             P@       Q      X                   �?F�4�Dj�?&            �M@        R      U                   �?�q�q�?             .@        S      T                `�X!@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        V      W                    @      �?              @       ������������������������       �                     @        ������������������������       �                     �?        Y      d                �!B@��2(&�?             F@       Z      c                   �?�����?             E@       [      b                @3�@�KM�]�?             C@       \      ]                �?�@��s����?             5@       ������������������������       �                     0@        ^      _                  �A@z�G�z�?             @        ������������������������       �                     @        `      a                  �D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     1@        ������������������������       �                     @        ������������������������       �                      @        f      g                   �?���Q��?             @        ������������������������       �                     �?        h      i                `f�.@      �?             @        ������������������������       �                     �?        j      k                  �A@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h*h-K ��h/��R�(KMmKK��h]�B�       �{@      q@      *@      :@      @      8@      @      @               @      @       @      @                       @              4@      $@       @      @              @       @       @              �?       @      �?                       @     �z@     �n@     r@     �a@      <@     �B@      8@      9@      3@      5@      .@      @      @              $@      @      @      @               @      @      @      @                      @      @              @      ,@              &@      @      @      �?      @              @      �?              @              @      @              @      @      �?       @              @      �?      @                      �?      @      (@       @      &@       @       @      �?      �?      �?                      �?      �?      @              @      �?       @               @      �?                      @       @      �?      �?      �?              �?      �?              �?             Pp@     �Y@     Pp@     �X@      e@      H@      3@      *@       @      @              @       @              1@      "@              �?      1@       @              @      1@       @      @       @      @       @       @              �?       @      @              &@             �b@     �A@     @P@      >@      "@              L@      >@      @      4@              @      @      1@      @      1@      @      ,@      �?              @      ,@       @              �?      ,@              �?      �?      *@      �?      &@              �?      �?      $@               @      �?      @               @      �?      �?      �?                      �?       @             �H@      $@      G@      "@      ;@      @      @       @       @              @       @               @      @              5@       @      @              1@       @      @      �?      @      �?      �?              (@      �?      @               @      �?      @      �?      @              3@      @      @              .@      @       @       @      �?              �?       @               @      �?              *@      @      &@      �?      @      �?      �?      �?      �?                      �?      @              @               @       @              �?       @      �?       @                      �?      @      �?       @              �?      �?              �?      �?             @U@      @      @       @              �?      @      �?       @      �?      @             �S@      @       @      �?      @      �?      �?      �?      �?                      �?      @               @             �Q@       @      �?             �Q@       @      @       @      @      �?      @      �?       @      �?      �?              @                      �?     �O@              W@     �I@     �P@     �I@      >@      *@              @      >@      "@      5@      @      2@      �?      &@              @      �?              �?      @              @      @       @              �?      @      �?      �?              �?      �?                       @      "@      @              @      "@       @      �?      �?              �?      �?               @      �?      @      �?      @              �?      �?              �?      �?              @              B@      C@       @      &@      �?      "@      �?                      "@      �?       @               @      �?              A@      ;@     �@@      6@      3@      @              @      3@      �?       @      �?              �?       @              &@              ,@      2@               @      ,@      $@       @      "@               @       @      @       @                      @      (@      �?      @      �?      @              �?      �?      �?                      �?      @              �?      @               @      �?      @              �?      �?       @      :@                      @     @a@     �Z@     �Q@      V@     �P@     �P@      E@      I@      C@      I@     �A@      B@      7@      2@              *@      7@      @      $@       @      @              @       @      @       @      �?              *@      @      @               @      @      @      @      @      @      @       @       @       @       @                      �?      @              �?              (@      2@              *@      (@      @      &@      @      @      @      �?               @      @               @       @       @       @                       @       @      �?       @      �?       @                      �?      @              �?              @      ,@              "@      @      @              @      @              @              9@      1@              (@      9@      @      ,@      @      (@      @      @      @      @      �?              �?      @               @       @              �?       @      �?              �?       @              @               @      �?      �?              �?      �?              �?      �?              &@      �?      @      �?      @                      �?      @              @      5@              .@      @      @      @      @               @      @       @      @                       @               @      Q@      2@      @      @              �?      @      @              @      @              O@      *@     �K@      *@      @             �I@      *@      H@      &@      $@      @      @      @      @                      @      @      �?      @                      �?      C@      @      C@      @      A@      @      1@      @      0@              �?      @              @      �?      �?      �?                      �?      1@              @                       @      @       @      �?               @       @      �?              �?       @               @      �?              @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ��~hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM=huh*h-K ��h/��R�(KM=��h|�B@O                         ��gS@l��n�?�           @�@              m                 `f�$@�xt��?�           ��@                                   /@.�ȓ�<�?�            �o@        ������������������������       �                     @                                  �4@�\��z�?�            `o@                                   �?`Ӹ����?            �F@        ������������������������       �                     @                                   �?�7��?            �C@        	       
                    3@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     B@                                    @(���g��?�            �i@        ������������������������       �                     @               *                    �?rLTAf�?}            �h@               !                    @k��9�?            �F@                               ���@�n`���?             ?@                                   �?$�q-�?             *@                                ���@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                                   �?�E��ӭ�?             2@                               �&B@"pc�
�?             &@                                  �?�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @                                    �?և���X�?             @                               �&B@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        "       #                    �?@4և���?             ,@        ������������������������       �                     @        $       %                   #@�C��2(�?             &@        ������������������������       �                     @        &       )                    �?z�G�z�?             @       '       (                    I@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        +       <                   �;@T����?f            @c@        ,       -                 ��@R���Q�?             D@        ������������������������       �                     @        .       9                    �?4?,R��?             B@       /       8                   �:@<���D�?            �@@       0       7                   �5@`Jj��?             ?@        1       2                    �?؇���X�?	             ,@        ������������������������       �                     �?        3       6                 �1@8�Z$���?             *@        4       5                  s@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     1@        ������������������������       �                      @        :       ;                   �9@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        =       j                 ���"@x�}b~|�?K            �\@       >       S                    �?��X��?I             \@        ?       F                  s�@$G$n��?            �B@       @       A                 ���@���N8�?             5@        ������������������������       �                     "@        B       E                    �?�8��8��?             (@       C       D                   @<@      �?              @       ������������������������       �z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     @        G       R                 �� @      �?             0@       H       K                    �?����X�?
             ,@        I       J                   �<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        L       Q                 ��(@      �?             (@       M       N                   �<@���!pc�?             &@       ������������������������       �؇���X�?             @        O       P                    >@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        T       i                    �?Х-��ٹ?1            �R@       U       \                 �?�@@-�_ .�?0            �R@        V       W                 ���@ ���J��?            �C@        ������������������������       �        
             1@        X       [                 �&B@���7�?             6@        Y       Z                   �=@z�G�z�?             @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �        
             1@        ]       h                    �?�#-���?            �A@       ^       a                 @3�@�C��2(�?            �@@        _       `                   �D@���Q��?             @       ������������������������       �      �?             @        ������������������������       �                     �?        b       g                 ��i @h�����?             <@       c       d                    ?@���N8�?             5@        ������������������������       �                     (@        e       f                   �@@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        k       l                    ?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        n                          @r�qu�?�             x@       o       �                  x#J@B��C���?�            u@       p       �                 `f�C@~�����?�            `r@       q       �                   �A@��(%��?�            Pq@       r       �                   �>@S9����?�            �p@       s       �                    �?     ��?�             p@       t       �                    �?�0{9��?u            �g@        u       v                 P�>,@Ԫ2��?%            �L@        ������������������������       �                     9@        w       �                    �?      �?             @@       x       y                 pF�-@��a�n`�?             ?@        ������������������������       �                      @        z       �                   �H@д>��C�?             =@       {       �                   �6@ȵHPS!�?             :@        |       }                     @���!pc�?             &@        ������������������������       �                     �?        ~       �                    ;@z�G�z�?             $@               �                 @3�/@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     .@        �       �                     �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                     �?��ׂ�?P            ``@        �       �                   @>@��+��?            �B@       �       �                    �?`՟�G��?             ?@        �       �                 �ܵ<@      �?              @        ������������������������       �                     @        �       �                   �E@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                 03k:@\X��t�?             7@        �       �                   �?@�q�q�?             @        ������������������������       �                     �?        �       �                   �9@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 `f�;@ҳ�wY;�?             1@       �       �                   �J@�q�q�?	             (@       �       �                   @B@r�q��?             @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     @        �       �                   @=@z�G�z�?             @        ������������������������       �                     �?        �       �                   @K@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �J@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?��8��)�?9            �W@        �       �                 @Q,@�	j*D�?             *@        ������������������������       �                     �?        �       �                     @      �?             (@        ������������������������       �                     @        �       �                    �?���Q��?             @       �       �                 `v�0@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?xdQ�m��?2            @T@       �       �                   @N@���N8�?&            �O@       �       �                     @�]0��<�?$            �N@       �       �                 `fF)@`�q�0ܴ?            �G@        ������������������������       �        	             2@        �       �                   �*@ 	��p�?             =@       �       �                    @@�����?             5@       ������������������������       �                     .@        �       �                    G@�q�q�?             @       �       �                    C@      �?             @        ������������������������       �      �?              @        ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     ,@        �       �                   �P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                     @�����H�?             2@       �       �                   �@@؇���X�?	             ,@        �       �                   �7@�q�q�?             @        ������������������������       �                     @        �       �                   �<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �*@.Lj���?0             Q@        ������������������������       �                     $@        �       �                    #@>n�T��?+             M@        ������������������������       �        
             *@        �       �                    �?�ݏ^���?!            �F@       �       �                    ,@�q�q�?            �@@        ������������������������       �                      @        �       �                 pF�,@¦	^_�?             ?@        ������������������������       �                      @        �       �                    �?>���Rp�?             =@       �       �                   �:@������?             ;@        ������������������������       �                      @        �       �                    �?p�ݯ��?             3@        ������������������������       �                     "@        �       �                   �H@�z�G��?             $@       �       �                 `v�5@�<ݚ�?             "@        ������������������������       �                      @        �       �                    �?����X�?             @        ������������������������       �                     �?        �       �                    @r�q��?             @       �       �                 ���9@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     (@        ������������������������       �                     $@        �       �                   B@���!pc�?             &@        ������������������������       �                      @        �       �                    �?�q�q�?             "@       �       �                    �?      �?             @       �       �                 �DpB@      �?             @        �       �                    +@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?������?             1@        �       �                    �?���Q��?             @       �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    H@�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        �                       �R@8�$�>�?            �E@       �                         �G@������?             A@       �                          �?؇���X�?             <@       �       �                    �?z�G�z�?             4@        ������������������������       �                     @        �                          >@�	j*D�?             *@        �                            @z�G�z�?             @                              ���M@      �?             @                                7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @              	                   �?�q�q�?             @        ������������������������       �                      @        
                         O@      �?             @        ������������������������       �                      @        ������������������������       �                      @                                 �?�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @                                 @�*/�8V�?            �G@                                =@r�q��?             >@                             ��T?@�>����?             ;@       ������������������������       �                     5@                                 �?�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     1@              .                   �?�MI8d�?-            �R@             '                pf�Z@D>�Q�?             J@             "                   �?<���D�?            �@@                                 �?d}h���?	             ,@       ������������������������       �                      @                              ��hU@      �?             @        ������������������������       �                      @               !                   �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        #      $                   �?�}�+r��?             3@       ������������������������       �        	             0@        %      &                03U@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        (      )                ���[@�d�����?             3@        ������������������������       �                      @        *      +                 "�`@@�0�!��?
             1@        ������������������������       �                     @        ,      -                   �?���!pc�?             &@       ������������������������       �                      @        ������������������������       �                     @        /      <                  �m@��2(&�?             6@       0      ;                `fmj@d}h���?
             ,@       1      2                   �?8�Z$���?	             *@        ������������������������       �                     @        3      8                ���`@�q�q�?             @       4      7                ���X@      �?             @       5      6                  �F@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        9      :                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �t�b�`     h�h*h-K ��h/��R�(KM=KK��h]�B�       {@     pq@     Pz@      k@     �i@      I@              @     �i@     �G@     �E@       @      @             �B@       @      �?       @               @      �?              B@              d@     �F@      @             @c@     �F@      3@      :@      @      9@      �?      (@      �?      @      �?                      @              @      @      *@       @      "@       @      @              @       @                       @      @      @       @      @       @                      @      �?              *@      �?      @              $@      �?      @              @      �?       @      �?       @                      �?       @             �`@      3@      ?@      "@              @      ?@      @      =@      @      =@       @      (@       @      �?              &@       @      @       @      @                       @       @              1@                       @       @      �?              �?       @              Z@      $@     �Y@      "@      @@      @      4@      �?      "@              &@      �?      @      �?      @      �?      @              @              (@      @      $@      @      �?      �?      �?                      �?      "@      @       @      @      @      �?       @       @               @       @              �?               @             �Q@      @     �Q@      @      C@      �?      1@              5@      �?      @      �?      �?      �?      @              1@              @@      @      >@      @      @       @      @      �?              �?      ;@      �?      4@      �?      (@               @      �?              �?       @              @               @              �?              �?      �?              �?      �?              k@     �d@     �e@     @d@      d@     �`@     `b@     @`@      b@     �^@     �`@     �^@     �[@     @S@       @     �H@              9@       @      8@      @      8@       @              @      8@      @      7@      @       @      �?               @       @       @      �?              �?       @                      @              .@       @      �?       @                      �?      �?             �Y@      <@      2@      3@      1@      ,@      @      @      @              �?      @              @      �?              *@      $@       @      @      �?              �?      @      �?                      @      &@      @      @      @      �?      @      �?      �?              @      @              @      �?      �?              @      �?      @                      �?      �?      @              @      �?             @U@      "@      "@      @              �?      "@      @      @               @      @      �?      @      �?                      @      �?              S@      @      N@      @     �M@       @     �F@       @      2@              ;@       @      3@       @      .@              @       @       @       @      �?      �?      �?      �?       @               @              ,@              �?      �?              �?      �?              0@       @      (@       @      @       @      @              �?       @      �?                       @       @              @              7@     �F@              $@      7@     �A@              *@      7@      6@      &@      6@       @              "@      6@       @              @      6@      @      4@               @      @      (@              "@      @      @      @       @       @              @       @              �?      @      �?      @      �?      @                      �?       @                      �?               @      (@              $@              @       @               @      @      @      @      @      @      �?      �?      �?              �?      �?               @                       @              @      *@      @       @      @       @      �?              �?       @                       @      &@      �?      &@                      �?      .@      <@       @      :@      @      8@      @      0@              @      @      "@      @      �?      @      �?      �?      �?      �?                      �?       @              �?                       @               @      @       @       @               @       @               @       @              @       @               @      @              E@      @      9@      @      9@       @      5@              @       @      @                       @              @      1@              (@      O@      "@     �E@      @      =@      @      &@               @      @      @       @              �?      @              @      �?              �?      2@              0@      �?       @      �?                       @      @      ,@       @              @      ,@              @      @       @               @      @              @      3@      @      &@       @      &@              @       @      @      �?      @      �?       @               @      �?                      �?      �?      �?      �?                      �?      �?                       @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ��.hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM!huh*h-K ��h/��R�(KM!��h|�B@H         t                     @<��z��?�           @�@               	                    .@
;&����?�             t@                                    �?�����H�?             ;@                                   @      �?              @                                   �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        	             3@        
       %                    �?,K/c��?�            pr@                                   �?">�֕�?.            �Q@        ������������������������       �                     >@               $                     �?�G�z��?             D@              !                    �?�P�*�?             ?@                               `f�B@�f7�z�?             =@                                �ܵ<@"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@                                   �?X�<ݚ�?             2@                               p�w@���|���?	             &@                                  �?�z�G��?             $@       ������������������������       �                     @                                  �5@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?                                Ȉ�Q@և���X�?             @        ������������������������       �                     �?                                   @K@�q�q�?             @                               �̾w@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        "       #                    6@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        &       9                    �?v�(��O�?�             l@        '       0                     �?`<)�+�?8            @S@        (       )                    �?@-�_ .�?            �B@       ������������������������       �                     ;@        *       +                    �?z�G�z�?             $@        ������������������������       �                     @        ,       -                   �8@�q�q�?             @        ������������������������       �                     @        .       /                 ���`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        1       8                    �?�(\����?!             D@       2       7                   �*@h�����?             <@       3       6                   �9@@4և���?             ,@        4       5                   �6@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �        
             &@        ������������������������       �                     ,@        ������������������������       �        	             (@        :       W                     �?�x
�2�?_            �b@        ;       V                    R@d��0u��?(             N@       <       =                 ��$:@$gv&��?'            �M@        ������������������������       �                     *@        >       ?                    �?��+7��?!             G@        ������������������������       �                     �?        @       S                   �E@������?             �F@       A       L                    �?���Q��?             9@       B       K                    �?ҳ�wY;�?             1@       C       J                   �@@���Q��?             .@       D       I                   �>@"pc�
�?	             &@        E       F                 `fF<@���Q��?             @        ������������������������       �      �?              @        G       H                   �<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        M       P                 `f�N@      �?              @        N       O                    9@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        Q       R                 03U@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        T       U                    �?ףp=
�?             4@       ������������������������       �                     2@        ������������������������       �                      @        ������������������������       �                     �?        X       s                    �?h�V���?7             V@       Y       d                    &@������?*            �Q@        Z       [                    @�d�����?             3@        ������������������������       �                     @        \       a                   �H@X�Cc�?             ,@       ]       `                   �5@�<ݚ�?             "@        ^       _                   �1@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     @        b       c                   �P@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        e       f                    �?�:�]��?            �I@        ������������������������       �                     �?        g       r                    �?HP�s��?             I@       h       i                   �;@dP-���?            �G@        ������������������������       �                     8@        j       q                   @A@�㙢�c�?             7@        k       n                    =@      �?              @        l       m                   �*@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        o       p                    @@���Q��?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �        	             .@        ������������������������       �                     @        ������������������������       �                     2@        u       �                    �?r9��X��?�            `x@        v       �                 ��Y7@���Q��?I             ^@       w       x                    �?`Y���?9            �V@        ������������������������       �                     @        y       �                 �̌@d�
��?6             V@        z       {                    �?l��
I��?             ;@        ������������������������       �                     @        |       }                   �3@�ՙ/�?             5@        ������������������������       �                     @        ~                        ���@������?             1@        ������������������������       �                     @        �       �                 �Y5@���|���?	             &@       �       �                    �?X�<ݚ�?             "@       �       �                    9@      �?              @        ������������������������       �                     �?        �       �                    �?և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ��.@��7��?$            �N@       �       �                    �?R���Q�?             D@        �       �                 P��+@�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        �       �                    3@�n`���?             ?@        �       �                    $@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?ȵHPS!�?             :@       �       �                 ���#@     ��?	             0@       �       �                   �9@@4և���?             ,@        ������������������������       �                     "@        �       �                   �;@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     $@        �       �                    ;@�q�q�?             5@        �       �                    �?����X�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �?؇���X�?             ,@        ������������������������       �                      @        ������������������������       �                     (@        �       �                 ��T?@ܷ��?��?             =@       ������������������������       �        	             2@        �       �                 ��p@@���!pc�?             &@        ������������������������       �                     @        ������������������������       �                      @        �                           �?l ��H|�?�            �p@       �       �                 �� @Ί�C�o�?�            �o@        ������������������������       �                     @        �       �                   �0@� ��?�             o@        �       �                     @�q�q�?             8@       �       �                    �?և���X�?	             ,@       �       �                    &@      �?              @        ������������������������       �                     �?        �       �                 pf�@����X�?             @        ������������������������       �                      @        �       �                 �̌!@���Q��?             @       ������������������������       �      �?             @        ������������������������       �                     �?        �       �                    ,@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        �                          �?�r����?�             l@       �       �                    �?�I�,ѽ�?�            @g@        �       �                    ;@d}h���?             <@        �       �                 ��y@և���X�?             @        ������������������������       �                     �?        �       �                 xF*@�q�q�?             @       �       �                    5@���Q��?             @        ������������������������       �                      @        �       �                   �7@�q�q�?             @       �       �                 ���@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ���@�����?             5@        ������������������������       �                      @        �       �                    ?@8�Z$���?             *@       �       �                   �<@z�G�z�?	             $@       �       �                   @<@�����H�?             "@       �       �                   @@      �?              @       ������������������������       �r�q��?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �>@���1���?n            �c@       �       �                   �;@���^���?P            �\@       �       �                   �:@ܷ��?��?-             M@       �       �                 �!&B@x�}b~|�?,            �L@       �       �                 ��L@@4և���?+             L@        �       �                    �?R���Q�?             4@        ������������������������       �                     @        �       �                   �4@@�0�!��?             1@        ������������������������       �                     @        �       �                 �?$@�θ�?	             *@       �       �                 ���@�����H�?             "@        �       �                 �&b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �6@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �3@������?             B@        �       �                 ��Y @@4և���?
             ,@        �       �                 �?�@      �?             @        ������������������������       �                      @        ������������������������       �      �?              @        ������������������������       �                     $@        ������������������������       �                     6@        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   @<@���U�?#            �L@       �       �                  sW@`2U0*��?             I@        �       �                    �?�C��2(�?             &@       ������������������������       �                     @        �       �                 pf�@r�q��?             @        ������������������������       �                      @        ������������������������       �      �?             @        �       �                 ��) @ ���J��?            �C@       ������������������������       �                     ;@        �       �                 pf� @�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     @        �       �                 �&B@RB)��.�?            �E@        ������������������������       �                     3@        �       �                   �@      �?             8@        ������������������������       �                      @        �                         @@@�X����?             6@        �       �                 �?�@      �?              @        ������������������������       �                     �?                                 �?@����X�?             @        ������������������������       �                     �?                              d�6@@�q�q�?             @                             ��i @���Q��?             @                             @3�@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        	                      @3�@؇���X�?
             ,@        
                      �?�@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @                                 �?:�&���?            �C@                                �?�θ�?             :@                                �?���N8�?             5@        ������������������������       �                     @                              ��@�E��ӭ�?             2@        ������������������������       �                     @                              pf�'@�q�q�?             (@                                �9@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @                                 �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @                               �v6@$�q-�?             *@       ������������������������       �                     "@                              03�7@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             2@        �t�bh�h*h-K ��h/��R�(KM!KK��h]�B       p|@     p@     @c@      e@      @      8@      @      @      @       @      @                       @              @              3@     �b@      b@      6@      H@              >@      6@      2@      *@      2@      (@      1@       @      "@       @                      "@      $@       @      @      @      @      @      @              �?      @      �?                      @              �?      @      @      �?               @      @       @      �?       @                      �?              @      �?      �?              �?      �?              "@              `@      X@      @     �R@       @     �A@              ;@       @       @              @       @      @              @       @      �?              �?       @              �?     �C@      �?      ;@      �?      *@      �?       @              �?      �?      �?              &@              ,@              (@     �_@      6@     �G@      *@     �G@      (@      *@              A@      (@      �?             �@@      (@      .@      $@      &@      @      "@      @      "@       @      @       @      �?      �?       @      �?              �?       @              @                      @       @              @      @      �?      @      �?                      @      @      �?      @                      �?      2@       @      2@                       @              �?     �S@      "@     �N@      "@      ,@      @      @              "@      @      @       @       @       @      �?              �?       @      @               @      @              @       @             �G@      @      �?              G@      @     �E@      @      8@              3@      @      @      @      �?       @               @      �?              @       @       @              �?       @      .@              @              2@             �r@     @V@      R@      H@      G@     �F@              @      G@      E@       @      3@              @       @      *@      @              @      *@              @      @      @      @      @      @      @              �?      @      @              @      @              �?                       @      C@      7@      ?@      "@      @      @              @      @              9@      @       @      @       @                      @      7@      @      *@      @      *@      �?      "@              @      �?              �?      @                       @      $@              @      ,@      @       @      @                       @       @      (@       @                      (@      :@      @      2@               @      @              @       @             �l@     �D@     `j@     �D@              @     `j@      C@      0@       @      @       @      @      @              �?      @       @       @              @       @       @       @      �?              �?      @              @      �?              $@             `h@      >@     `d@      7@      6@      @      @      @      �?               @      @       @      @               @       @      �?      �?      �?              �?      �?              �?                      �?      3@       @       @              &@       @       @       @       @      �?      @      �?      @      �?       @              �?                      �?      @             �a@      1@     �Z@       @      J@      @      J@      @      J@      @      1@      @      @              ,@      @      @              $@      @       @      �?      �?      �?      �?                      �?      @               @       @               @       @             �A@      �?      *@      �?      @      �?       @              �?      �?      $@              6@                      �?              �?     �K@       @      H@       @      $@      �?      @              @      �?       @              @      �?      C@      �?      ;@              &@      �?              �?      &@              @              A@      "@      3@              .@      "@               @      .@      @      @      @      �?               @      @              �?       @      @       @      @      �?      @      �?       @              �?      �?                      �?      (@       @      @       @      @                       @       @              @@      @      4@      @      0@      @      @              *@      @      @              @      @      �?      @              @      �?              @              @      �?              �?      @              (@      �?      "@              @      �?              �?      @              2@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�DhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B�@         �                    �?��6���?�           @�@              ;                    �?2�E���?Y           ��@                                    @�������?g            `d@                                   �?      �?<             X@       ������������������������       �        "             K@                                   �?@4և���?             E@        ������������������������       �                     @                                  �7@�#-���?            �A@       	                          �;@�����H�?             ;@        
                          �9@���Q��?             @        ������������������������       �                     �?                                   �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     6@        ������������������������       �                      @                                   �?�萻/#�?+            �P@                                  �+@      �?              @        ������������������������       �                     �?                                �%@����X�?             @        ������������������������       �                      @        ������������������������       �                     @                                  �4@Ɣ��Hr�?%            �M@                                �L�@���!pc�?             &@        ������������������������       �                     @                                   �?      �?             @        ������������������������       �                      @                                   3@      �?             @        ������������������������       �                     �?        ������������������������       �                     @               (                 �̌@     ��?             H@                !                    ;@HP�s��?             9@        ������������������������       �                     &@        "       #                 ���@؇���X�?	             ,@        ������������������������       �                     �?        $       %                 ���@$�q-�?             *@        ������������������������       �                     @        &       '                 �&B@�����H�?             "@       ������������������������       �؇���X�?             @        ������������������������       �                      @        )       2                   p"@\X��t�?             7@        *       +                    �?ףp=
�?             $@        ������������������������       �                     �?        ,       -                    :@�����H�?             "@        ������������������������       �                     @        .       1                 @3�@z�G�z�?             @        /       0                 �?�@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        3       4                    �?�	j*D�?             *@        ������������������������       �                     �?        5       :                    @@�q�q�?             (@       6       7                    ;@�q�q�?             @        ������������������������       �                      @        8       9                 ��1@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        <       �                 ��$:@s�As��?�            w@       =       �                    �?�)���Y�?�            `r@       >       Q                 ��@�'��?�            �q@        ?       P                    �?`Ql�R�?9            �W@       @       A                     @�d���?6            �U@        ������������������������       �                     "@        B       I                    �? ���J��?1            �S@        C       H                 ���@ �q�q�?             8@       D       E                 03S@      �?	             0@        ������������������������       �                     @        F       G                   �7@�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                      @        J       K                    �?@3����?"             K@        ������������������������       �                     4@        L       O                   �;@г�wY;�?             A@        M       N                    :@�IєX�?	             1@       ������������������������       �                     0@        ������������������������       �                     �?        ������������������������       �                     1@        ������������������������       �                     @        R       �                    �?�YM_b�?|            �g@       S       �                   @@@��D<j�?o            �e@       T                           ?@�����?R            �`@       U       ^                   @@��7PB��?M            �_@        V       Y                 �?$@      �?             ,@        W       X                    ;@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        Z       ]                   �9@X�<ݚ�?             "@       [       \                   �5@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        _       `                 @3�@�=|+g��?F            @\@        ������������������������       �                     9@        a       f                    �?�Ra����?7             V@        b       e                     @�q�q�?             @       c       d                 `��,@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        g       r                     @�̨�`<�?4            @U@        h       k                    &@PN��T'�?             ;@        i       j                   �6@�<ݚ�?             "@        ������������������������       ��q�q�?             @        ������������������������       �                     @        l       m                   �;@�����H�?             2@       ������������������������       �        	             ,@        n       q                    =@      �?             @       o       p                   �*@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        s       z                 ��i @��ϭ�*�?#             M@        t       u                   �1@PN��T'�?             ;@        ������������������������       �                     �?        v       w                   �3@ȵHPS!�?             :@        ������������������������       ��q�q�?             @        x       y                 ��) @���}<S�?             7@       ������������������������       �                     5@        ������������������������       �                      @        {       |                   �<@�g�y��?             ?@       ������������������������       �                     <@        }       ~                 ���"@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 ��i @և���X�?             @       �       �                   �@z�G�z�?             @        ������������������������       �                      @        �       �                 �?�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                     @ ���J��?            �C@        �       �                 ��Y)@�8��8��?             (@        ������������������������       �                     @        �       �                   �*@      �?              @        �       �                    E@      �?             @       ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     ;@        �       �                    �?     ��?             0@        ������������������������       �                      @        �       �                   �4@d}h���?             ,@        ������������������������       �                      @        �       �                     @�8��8��?
             (@        ������������������������       �                     @        �       �                 �&B@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        �       �                   �8@�O�y���?7            �R@        ������������������������       �                     @        �       �                   �;@ꮃG��?2            @Q@        ������������������������       �                     &@        �       �                    �?>n�T��?,             M@       �       �                   �L@�+��<��?!            �E@       �       �                   �G@Hث3���?            �C@       �       �                   �F@     ��?             @@       �       �                    �?l��[B��?             =@        �       �                 ���<@�q�q�?             "@        ������������������������       �                     @        �       �                   �A@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                      @�G�z��?             4@       �       �                   �>@      �?             0@        �       �                   �E@�����H�?             "@       ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     @        �       �                    >@      �?             @        ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �J@����X�?             @        ������������������������       �                     @        �       �                   �K@�q�q�?             @        ������������������������       �                     �?        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                     �?������?             .@       �       �                 03�M@���Q��?             $@        ������������������������       �                     �?        �       �                   �G@�q�q�?             "@       ������������������������       �                     @        �       �                 @�pX@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ���S@����E��?i            �f@       �       �                    @B�F<��?Z             c@       �       �                    @r�J���?W            �b@       �       �                    #@�Jl$G��?A            �[@        �       �                     @�IєX�?             A@        ������������������������       �                     *@        �       �                    �?�����?             5@        �       �                    �?"pc�
�?             &@        ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                      @        �       �                   �&@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     $@        �       �                     @�eP*L��?/            @S@       �       �                    �?X�<ݚ�?            �F@       ������������������������       �                     9@        ������������������������       �        	             4@        �       �                    �?     ��?             @@       �       �                    �?      �?             2@        �       �                 03�-@X�<ݚ�?             "@        ������������������������       �                     @        �       �                    �?z�G�z�?             @        ������������������������       �                      @        �       �                   �<@�q�q�?             @       �       �                  S�2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �;@X�<ݚ�?             "@       �       �                    �?����X�?             @       �       �                    �?r�q��?             @        ������������������������       �                      @        �       �                 ��l4@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?@4և���?	             ,@        �       �                 ��&@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     (@        �       �                    �?�MI8d�?            �B@        ������������������������       �                     &@        �       �                   �6@�θ�?             :@       �       �                   �0@ҳ�wY;�?
             1@       �       �                    �?�8��8��?	             (@        ������������������������       �                     @        �       �                    @؇���X�?             @        �       �                     @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     @        �                          O@ �Cc}�?             <@       �       �                   kp@ ��WV�?             :@       ������������������������       �                     6@                                  5@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �t�bh�h*h-K ��h/��R�(KMKK��h]�B0       Pz@     0r@     0u@      h@      ?@     �`@      @     @W@              K@      @     �C@              @      @      @@      @      8@      @       @      �?               @       @               @       @                      6@               @      <@     �C@      @      @              �?      @       @               @      @              7@      B@       @      @      @              @      @               @      @      �?              �?      @              .@     �@@       @      7@              &@       @      (@      �?              �?      (@              @      �?       @      �?      @               @      *@      $@      "@      �?      �?               @      �?      @              @      �?      �?      �?      �?                      �?      @              @      "@              �?      @       @      @       @       @               @       @               @       @                      @     @s@     �N@     �p@      ;@      p@      ;@      W@       @     @U@       @      "@              S@       @      7@      �?      .@      �?      @              &@      �?              �?      &@               @             �J@      �?      4@             �@@      �?      0@      �?      0@                      �?      1@              @             �d@      9@     �b@      6@     @\@      5@     �[@      1@      @      @      @       @      @                       @      @      @      @       @               @      @                      @     �Y@      $@      9@             �S@      $@       @      �?      �?      �?              �?      �?              �?              S@      "@      7@      @      @       @      �?       @      @              0@       @      ,@               @       @      �?       @               @      �?              �?             �J@      @      7@      @              �?      7@      @       @      �?      5@       @      5@                       @      >@      �?      <@               @      �?       @                      �?      @      @      �?      @               @      �?       @      �?                       @       @              C@      �?      &@      �?      @              @      �?      @      �?      �?      �?       @              @              ;@              *@      @       @              &@      @               @      &@      �?      @              @      �?              �?      @              &@             �D@      A@      @             �A@      A@              &@     �A@      7@      8@      3@      4@      3@      2@      ,@      .@      ,@      @      @      @               @      @              @       @              "@      &@       @       @      �?       @              @      �?      �?      @              �?      @      �?      �?               @      @               @      @              @       @      �?      �?              �?      �?              �?      �?              @              &@      @      @      @              �?      @      @      @              �?      @              @      �?              @             �T@     �X@     �S@     @R@     �R@     @R@      F@     �P@       @      @@              *@       @      3@       @      "@              @       @      @               @       @      @       @                      @              $@      E@     �A@      4@      9@              9@      4@              6@      $@      "@      "@      @      @      @              �?      @               @      �?       @      �?      �?      �?                      �?              �?      @      @       @      @      �?      @               @      �?      @              @      �?              �?               @              *@      �?      �?      �?      �?                      �?      (@              ?@      @      &@              4@      @      &@      @      &@      �?      @              @      �?      �?      �?      �?                      �?      @                      @      "@              @              @      9@      �?      9@              6@      �?      @      �?                      @       @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ���MhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMShuh*h-K ��h/��R�(KMS��h|�B�T         ~                     @�U��h��?�           @�@               W                    �?�n�q�Z�?�            `s@              D                   �J@�҇���?�            �g@              C                   @M@6�;�vv�?f            @b@                                  �?��c:�?`            @a@                                   �?X�<ݚ�?             2@                                  �?��.k���?             1@               	                 `v7<@؇���X�?             @       ������������������������       �                     @        
                        hލC@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   �?�z�G��?	             $@                                 �L@�q�q�?             "@                                 @G@      �?              @                               ���<@����X�?             @        ������������������������       �                     @                                   �?      �?             @                                  A@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?                                   �?*;L]n�?P             ^@        ������������������������       �                    �A@               $                   �:@�����	�?:            @U@               #                    5@�}�+r��?             3@                                   �2@ףp=
�?             $@       ������������������������       �                      @        !       "                   �'@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        %       6                     �?r�q��?,            �P@        &       +                 `fF<@�������?             >@        '       (                 ��$:@��S�ۿ?
             .@       ������������������������       �                     $@        )       *                 03k:@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ,       -                   �;@���Q��?             .@        ������������������������       �                      @        .       5                   �J@�	j*D�?
             *@       /       4                   `@@�q�q�?	             (@        0       1                   �<@�q�q�?             @        ������������������������       �                     @        2       3                   @>@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        7       8                    @@�����H�?             B@        ������������������������       �        	             ,@        9       B                   �*@"pc�
�?             6@        :       A                   �F@�q�q�?             (@       ;       <                   �'@      �?              @        ������������������������       �                     �?        =       @                   @D@և���X�?             @       >       ?                   @B@���Q��?             @       ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                      @        E       R                    �?��s����?             E@       F       M                    �?z�G�z�?             9@       G       H                    �?      �?
             0@       ������������������������       �                     *@        I       J                  �}S@�q�q�?             @        ������������������������       �                     �?        K       L                   @D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        N       O                    �?X�<ݚ�?             "@        ������������������������       �                     @        P       Q                   �4@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        S       V                 ��gS@@�0�!��?             1@        T       U                 03�P@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     &@        X       u                 Ј�U@�̚��?L            �^@       Y       `                    �?J`mL�#�?<            @X@       Z       _                    �?p���?              I@       [       ^                   �6@`���i��?             F@        \       ]                 ��m1@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     E@        ������������������������       �                     @        a       d                   �3@p�v>��?            �G@        b       c                    *@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        e       l                    �?��P���?            �D@        f       k                    �?      �?              @       g       j                 ���S@      �?             @       h       i                 ��`E@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        m       p                     �?"pc�
�?            �@@        n       o                    =@8�Z$���?             *@        ������������������������       �                      @        ������������������������       �                     &@        q       r                    �?z�G�z�?             4@        ������������������������       �                      @        s       t                    +@�q�q�?             (@        ������������������������       �                     @        ������������������������       �                      @        v       }                    4@HP�s��?             9@        w       x                    �?���Q��?             @        ������������������������       �                     �?        y       z                    �?      �?             @        ������������������������       �                     �?        {       |                     @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     4@               >                ��Y7@!��)��?�             y@       �       �                  �#@`� ��?�            pu@       �       �                    �?4�=ݍ�?�            �o@       �       �                   �0@��mo*�?�            �m@        �       �                    �?�	j*D�?	             *@       ������������������������       �                      @        �       �                 P��@z�G�z�?             @        ������������������������       �                      @        �       �                 pFD!@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ���@�b<�J�?�            �k@        �       �                   �@@ �o_��?B             Y@       �       �                   �3@H���I�?6            �S@        ������������������������       �                      @        �       �                    �?:%�[��?0            �Q@        �       �                    �?؇���X�?             5@       �       �                    �?$�q-�?	             *@        ������������������������       �                     @        �       �                 ���@ףp=
�?             $@        ������������������������       �                     @        �       �                 �&B@؇���X�?             @       ������������������������       �z�G�z�?             @        ������������������������       �                      @        �       �                 ���@      �?              @        ������������������������       �                      @        �       �                 �&B@�q�q�?             @       �       �                   �7@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?z�G�z�?"             I@        �       �                 ���@8�Z$���?             :@       �       �                 ���@      �?
             (@        ������������������������       �                      @        �       �                    5@�z�G��?             $@        ������������������������       �                     �?        �       �                    9@�<ݚ�?             "@        ������������������������       �                     �?        �       �                    =@      �?              @       ������������������������       �����X�?             @        ������������������������       �                     �?        �       �                  s�@@4և���?             ,@        ������������������������       �                     @        �       �                 ��(@�C��2(�?             &@       �       �                   �<@      �?              @       ������������������������       �                     @        �       �                    >@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 P�N@      �?             8@       �       �                   �;@��s����?             5@       �       �                   �:@������?
             .@       �       �                 �&b@d}h���?	             ,@        ������������������������       �                      @        �       �                 ���@      �?             (@        ������������������������       �                     �?        �       �                 �?$@"pc�
�?             &@        ������������������������       �                     @        �       �                 �1@����X�?             @       �       �                   �5@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    :@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     5@        �       �                    �?n�6�Է�?M            �^@        �       �                 �� @z�G�z�?             $@       �       �                    ?@�<ݚ�?             "@       �       �                   �<@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                 �?�@4Ky\�?G            @\@        ������������������������       �                     @@        �       �                   �:@.�	F�9�?4            @T@        �       �                 pf� @P�Lt�<�?             C@        �       �                   �3@@4և���?
             ,@        ������������������������       �                     �?        ������������������������       �        	             *@        ������������������������       �                     8@        �       �                 @3�@�lg����?            �E@        �       �                   �?@�<ݚ�?             "@        ������������������������       �                     @        �       �                   �A@���Q��?             @        ������������������������       ��q�q�?             @        ������������������������       �      �?              @        �       �                 @!@�������?             A@       �       �                    �?�KM�]�?             3@       �       �                    �?�t����?             1@        ������������������������       �                     �?        �       �                 ��) @      �?             0@       �       �                    ?@@4և���?             ,@       ������������������������       �                      @        �       �                   �@@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ��y @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �;@��S���?             .@        ������������������������       �                     @        �       �                 ��)"@���!pc�?             &@        ������������������������       �                     @        �       �                 `f#@և���X�?             @        �       �                   �<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    I@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                 �&B@�����H�?
             2@        �       �                   �7@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     &@        �                         �8@��9܂�?5            @V@        �                          �?      �?             @@       �                          .@�q�����?             9@       �                          �?X�Cc�?	             ,@       �                          @�q�q�?             "@       �                          �?      �?              @                                 @����X�?             @                               �&@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?                                 �?���Q��?             @        ������������������������       �                     �?        	      
                   �?      �?             @        ������������������������       �                      @                                 @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                 �?���|���?             &@                                 �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                              �yW(@      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @              +                   �?�q�q�?"            �L@              "                   �?�ՙ/�?             5@                                 �?      �?             @                               S�2@�q�q�?             @                               �<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?              !                   �?�q�q�?             @                                 ;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        #      *                   �?�q�q�?             .@       $      %                   �?X�Cc�?             ,@        ������������������������       �                     @        &      '                   �?ףp=
�?             $@       ������������������������       �                     @        (      )                 �v6@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ,      =                   C@<ݚ)�?             B@       -      <                  @A@f���M�?             ?@       .      ;                   �?�θ�?             :@        /      6                   �?�q�q�?             "@       0      1                   �?�q�q�?             @        ������������������������       �                     �?        2      5                ��1@���Q��?             @       3      4                   ;@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        7      8                   <@�q�q�?             @        ������������������������       �                     �?        9      :                   >@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     1@        ������������������������       �                     @        ������������������������       �                     @        ?      N                   ?@�^����?#            �M@       @      A                   �?`�q�0ܴ?            �G@        ������������������������       �                     ;@        B      C                   �?ףp=
�?             4@        ������������������������       �                     @        D      G                   @�r����?             .@        E      F                pf�C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        H      I                �T�I@$�q-�?
             *@        ������������������������       �                     @        J      M                   �?r�q��?             @        K      L                   ;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        O      R                   �?�q�q�?             (@        P      Q                  �A@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �t�b�      h�h*h-K ��h/��R�(KMSKK��h]�B0       �z@     �q@     �`@      f@     @X@     �V@     @V@     �L@     @T@     �L@       @      $@       @      "@      �?      @              @      �?      �?      �?                      �?      @      @      @      @      @      @      @       @      @               @       @      �?       @               @      �?              �?                      �?      �?              �?                      �?     @R@     �G@             �A@     @R@      (@      2@      �?      "@      �?       @              �?      �?              �?      �?              "@             �K@      &@      7@      @      ,@      �?      $@              @      �?              �?      @              "@      @               @      "@      @       @      @       @      @              @       @      �?       @                      �?      @              �?              @@      @      ,@              2@      @       @      @      @      @      �?              @      @      @       @      �?       @       @                       @      @              $@               @               @      A@      @      4@      �?      .@              *@      �?       @              �?      �?      �?              �?      �?              @      @              @      @      �?              �?      @              @      ,@      @      @              @      @                      &@      B@     �U@      A@     �O@      �?     �H@      �?     �E@      �?      �?              �?      �?                      E@              @     �@@      ,@      �?      @      �?                      @      @@      "@      @      @      @      @      �?      @      �?                      @       @               @              ;@      @      &@       @               @      &@              0@      @       @               @      @              @       @               @      7@       @      @              �?       @       @      �?              �?       @               @      �?                      4@     �r@      Z@     �n@     @X@     �h@      M@     �f@      L@      @      "@               @      @      �?       @               @      �?              �?       @              f@     �G@      R@      <@     �I@      <@       @             �E@      <@      @      2@      �?      (@              @      �?      "@              @      �?      @      �?      @               @       @      @               @       @      @       @       @               @       @                       @      D@      $@      6@      @      "@      @       @              @      @              �?      @       @      �?              @       @      @       @      �?              *@      �?      @              $@      �?      @      �?      @              @      �?              �?      @              @              2@      @      1@      @      &@      @      &@      @       @              "@      @              �?      "@       @      @              @       @      @       @               @      @               @                      �?      @              �?       @      �?                       @      5@              Z@      3@       @       @      @       @       @       @       @                       @      @              �?              X@      1@      @@              P@      1@     �B@      �?      *@      �?              �?      *@              8@              ;@      0@       @      @              @       @      @      �?       @      �?      �?      9@      "@      1@       @      .@       @      �?              ,@       @      *@      �?       @              @      �?              �?      @              �?      �?              �?      �?               @               @      @              @       @      @      @              @      @      �?       @      �?                       @      @      �?      @                      �?      0@       @      @       @      @                       @      &@              I@     �C@      (@      4@      (@      *@      @      "@      @      @       @      @       @      @       @       @       @                       @              @              �?      �?               @      @      �?              �?      @               @      �?      �?      �?                      �?      @      @       @      �?       @                      �?      @      @              @      @                      @      C@      3@      *@       @      @      @      �?       @      �?      �?      �?                      �?              �?       @      �?      �?      �?              �?      �?              �?              $@      @      "@      @              @      "@      �?      @              @      �?      @                      �?      �?              9@      &@      4@      &@      4@      @      @      @       @      @              �?       @      @      �?      @      �?                      @      �?              �?       @              �?      �?      �?      �?                      �?      1@                      @      @              J@      @     �F@       @      ;@              2@       @      @              *@       @      �?      �?              �?      �?              (@      �?      @              @      �?       @      �?              �?       @              @              @      @       @      @              @       @              @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ9M�hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM+huh*h-K ��h/��R�(KM+��h|�B�J         >                    �?���y�?�           @�@               %                  I>@�p ��?M            �^@                               P�>,@0�� ��?'            �O@                                  �?\�Uo��?             C@                                 �9@<=�,S��?            �A@                                   �?ףp=
�?             $@        ������������������������       �                     @                                   5@      �?             @       	       
                 �{@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @                                  �=@�J�4�?             9@                                 �<@������?             1@                               ���@@4և���?
             ,@        ������������������������       �                     @                                  @@�C��2(�?             &@                                  �?�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @                                ��}@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @               $                    �?�J�4�?             9@              #                    �?���}<S�?             7@                                  6@8�Z$���?             *@        ������������������������       �                     @               "                     @      �?              @               !                 ��4=@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                      @        &       9                     �?������?&             N@       '       (                    �?�E��ӭ�?"             K@       ������������������������       �                     ;@        )       2                    �?X�<ݚ�?             ;@       *       +                 `f�A@�q�q�?	             2@        ������������������������       �                     @        ,       -                   �3@z�G�z�?             .@        ������������������������       �                     �?        .       /                   �?@؇���X�?             ,@       ������������������������       �                     "@        0       1                 �;|r@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        3       8                 �U�X@�q�q�?             "@       4       5                   �:@؇���X�?             @        ������������������������       �                     @        6       7                 ���S@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        :       =                 pV�C@r�q��?             @        ;       <                    0@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ?       �                    �?�����2�?t           h�@        @       �                    �?Rh6��p�?x            �h@       A       R                    �? �o_��?[            �b@        B       Q                 ��|$@���!pc�?            �@@       C       D                    1@8�A�0��?             6@        ������������������������       �                     @        E       F                    4@�\��N��?	             3@        ������������������������       �                     �?        G       P                 pF @X�<ݚ�?             2@       H       I                    9@�θ�?             *@        ������������������������       �                     �?        J       K                 ���@      �?             (@        ������������������������       �                     �?        L       M                  s�@"pc�
�?             &@        ������������������������       �                     @        N       O                 �&B@����X�?             @       ������������������������       ����Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     &@        S       Z                    '@�(�Tw��?K            @]@        T       Y                 pf�0@����X�?             @       U       X                    �?      �?             @       V       W                   �&@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        [       h                     @^(��I�?F            �[@       \       ]                     �?����˵�?(            �M@        ������������������������       �                     :@        ^       g                   �;@�C��2(�?            �@@        _       f                    6@���!pc�?             &@        `       a                   �6@      �?             @        ������������������������       �                      @        b       e                    �?      �?             @       c       d                   �'@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     6@        i       �                    C@Np�����?            �I@       j       �                   @.@8�A�0��?             F@       k       �                    �?      �?             A@       l       }                   �;@��}*_��?             ;@       m       n                 pf�@����X�?             5@        ������������������������       �                      @        o       |                    �?�����?             3@       p       {                    9@      �?	             0@       q       z                   �6@��
ц��?             *@       r       y                 �[$@���|���?             &@       s       x                  �#@�z�G��?             $@       t       u                    4@և���X�?             @        ������������������������       �                      @        v       w                 �̜!@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ~                           =@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    ;@ףp=
�?             $@        �       �                    9@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�q�q��?             H@        �       �                   �4@      �?              @        �       �                 `f7@      �?             @        ������������������������       �                      @        �       �                     @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                 03�;@�z�G��?             D@        ������������������������       �                     @        �       �                 ���i@@�0�!��?             A@       �       �                    @      �?             @@       �       �                 ��T?@PN��T'�?             ;@        ������������������������       �                     "@        �       �                     @�<ݚ�?             2@        �       �                 ���`@      �?              @       ������������������������       �                     @        ������������������������       �                     @        �       �                    @ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     @        ������������������������       �                      @        �       �                     �?ހ�\���?�            px@        �       �                    �?���Q��?(             N@       �       �                    �?Ɣ��Hr�?'            �M@       �       �                   �>@�û��|�?             G@       �       �                   �9@�eP*L��?            �@@        ������������������������       �                     @        �       �                 03k:@�q�q�?             ;@        ������������������������       �                     @        �       �                   @=@�û��|�?             7@       �       �                 `f�;@��S���?             .@       �       �                    K@��
ц��?             *@       �       �                   @G@      �?              @       �       �                   @B@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                   �<@      �?              @        ������������������������       �                     @        �       �                   @D@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        
             *@        �       �                    D@�n_Y�K�?             *@        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �       *                   �?��@u�\�?�            �t@       �       #                0�H@�`�=	�?�            Ps@       �       "                   @`Pj���?�            �r@       �                         �B@���Y.�?�            �q@       �       �                    )@h�! &,�?�            `q@        ������������������������       �                     $@        �                         �N@�NJa&��?�            �p@       �       �                   �0@TY��&\�?�            �p@        �       �                 �̌"@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                     @�L���?�            0p@        �       �                   @B@l��\��?*             Q@       �       �                 `fF)@�t����?             �I@        �       �                    @�nkK�?             7@        ������������������������       �                     @        �       �                    &@      �?	             0@       �       �                   �6@ףp=
�?             $@        ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�>4և��?             <@       �       �                   �*@���B���?             :@       �       �                   �;@      �?             0@        ������������������������       �                     @        �       �                    =@���Q��?             $@        ������������������������       �                      @        �       �                    @@      �?              @        ������������������������       �                     @        ������������������������       ����Q��?             @        �       �                    >@ףp=
�?             $@        ������������������������       �                     @        �       �                   �7@z�G�z�?             @        ������������������������       �                     �?        �       �                   �@@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        
             1@        �                          �?��Y���?            �g@       �       �                   �8@��;M��?x            @f@        �       �                 @3�@@9G��?$            �H@        �       �                 �?�@$�q-�?             :@       �       �                 �?$@ �q�q�?             8@       ������������������������       �        	             *@        �       �                 ��L@�C��2(�?             &@        �       �                   �5@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   �4@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     7@        �       �                    �?�|K��2�?T             `@        �       �                   `3@�C��2(�?             6@       �       �                    �?�}�+r��?             3@       �       �                 03�@�X�<ݺ?             2@        ������������������������       �                     @        �       �                    >@@4և���?	             ,@       ������������������������       ��C��2(�?             &@        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �                          �?�ʠ����?F            �Z@       �                       @3�@�=C|F�?<            �U@        �                          �>@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                �;@ �Cc}�?:             U@                              pf� @�q�q�?             "@                               �:@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @                                �?@HP�s��?5            �R@        	                        �<@г�wY;�?             A@       
                       sW@XB���?             =@                              pf�@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     9@        ������������������������       �                     @                              @3�@,���i�?            �D@                               @@@��<b���?             7@                              P�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @                              �?�@R���Q�?             4@       ������������������������       �                     0@                                �D@      �?             @       ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �        
             2@        ������������������������       �        
             4@        ������������������������       �                     *@                                 Q@      �?             @        ������������������������       �                      @        ������������������������       �                      @               !                  �>@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        	             2@        $      )                ��?P@X�<ݚ�?             "@       %      (                   >@r�q��?             @       &      '                   ;@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     6@        �t�bh�h*h-K ��h/��R�(KM+KK��h]�B�       �|@      p@      N@     �O@      F@      3@      7@      .@      6@      *@      �?      "@              @      �?      @      �?      �?      �?                      �?               @      5@      @      *@      @      *@      �?      @              $@      �?       @      �?              �?       @               @                      @       @              �?       @      �?                       @      5@      @      5@       @      &@       @      @              @       @      @      �?      @                      �?              �?      $@                       @      0@      F@      .@     �C@              ;@      .@      (@      (@      @              @      (@      @              �?      (@       @      "@              @       @      @                       @      @      @      �?      @              @      �?       @               @      �?               @              �?      @      �?      @              @      �?                       @     �x@      h@     �Q@     �_@      E@      [@      "@      8@      "@      *@              @      "@      $@      �?               @      $@      @      $@              �?      @      "@      �?               @      "@              @       @      @       @      @               @      @                      &@     �@@      U@      @       @       @       @       @      �?       @                      �?              �?      @              <@     �T@      @      L@              :@      @      >@      @       @      @      @               @      @      �?      �?      �?              �?      �?               @                      @              6@      9@      :@      2@      :@      1@      1@      $@      1@      @      .@               @      @      *@      @      $@      @      @      @      @      @      @      @      @       @              �?      @              @      �?                      @      �?               @                      @              @      @       @      @                       @      @              �?      "@      �?      �?              �?      �?                       @      @              =@      3@      �?      @      �?      @               @      �?      �?              �?      �?                      @      <@      (@              @      <@      @      <@      @      7@      @      "@              ,@      @      @      @              @      @              "@      �?              �?      "@              @                       @     Pt@     �P@      B@      8@      B@      7@      <@      2@      .@      2@      @              "@      2@              @      "@      ,@       @      @      @      @      �?      @      �?      @              �?      �?      @              @      @               @              �?      @              @      �?       @      �?                       @      *@               @      @              @       @                      �?     r@      E@     �p@      E@     pp@     �B@     �n@     �B@     `n@     �A@              $@     `n@      9@      n@      7@      @       @               @      @             �m@      5@      O@      @     �F@      @      6@      �?      @              .@      �?      "@      �?      �?      �?       @              @              7@      @      5@      @      (@      @      @              @      @               @      @       @      @              @       @      "@      �?      @              @      �?      �?              @      �?              �?      @               @              1@              f@      .@     `d@      .@     �G@       @      8@       @      7@      �?      *@              $@      �?      @      �?              �?      @              @              �?      �?              �?      �?              7@              ]@      *@      4@       @      2@      �?      1@      �?      @              *@      �?      $@      �?      @              �?               @      �?       @                      �?      X@      &@      S@      &@      �?       @               @      �?             �R@      "@      @      @      @      �?      @                      �?               @     @Q@      @     �@@      �?      <@      �?      @      �?      �?               @      �?      9@              @              B@      @      2@      @      �?       @              �?      �?      �?      1@      @      0@              �?      @      �?      �?               @      2@              4@              *@               @       @               @       @               @       @               @       @              2@              @      @      �?      @      �?      @              �?      �?       @               @      @              6@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJpVhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B@G         \                    �?T�����?�           @�@                                   �?������?�             l@                                    @dP-���?            �G@       ������������������������       �                     A@               
                    �?�	j*D�?	             *@                               P��+@���|���?             &@        ������������������������       �                     @               	                 033.@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @               Q                   �=@PN���?s            @f@              H                    @�m��Wv�?I             [@              #                     @t]����?=            �V@                                   �?8�Z$���?            �C@        ������������������������       �                     �?                                 ���`@�S����?             C@                                   �?(N:!���?            �A@        ������������������������       �                      @                                  �9@PN��T'�?             ;@                                  �?�}�+r��?             3@                                   �?؇���X�?             @                                 �6@      �?             @        ������������������������       �                      @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     (@                                   �?      �?              @       ������������������������       �                     @                                  �7@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        !       "                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        $       C                    �?��B����?"             J@       %       8                   �:@      �?             G@       &       '                    �?���!pc�?             6@        ������������������������       �                     �?        (       7                    �?���N8�?             5@       )       *                    �?      �?             4@        ������������������������       �                      @        +       6                    �?�E��ӭ�?             2@       ,       -                 pf�@�eP*L��?             &@        ������������������������       �                      @        .       5                  �#@�q�q�?             "@       /       0                    4@؇���X�?             @        ������������������������       �                      @        1       4                   �6@z�G�z�?             @        2       3                 �̜!@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        9       B                   �<@�q�q�?             8@       :       A                    �?��+7��?             7@       ;       >                    �?�����?             3@       <       =                 pF @8�Z$���?             *@       ������������������������       �                     &@        ������������������������       �                      @        ?       @                    �?�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        D       G                    �?�q�q�?             @       E       F                 ��"@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        I       J                    �?@�0�!��?             1@        ������������������������       �                     @        K       L                      @�θ�?	             *@        ������������������������       �                      @        M       P                    @�C��2(�?             &@        N       O                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        R       [                    @������?*            �Q@       S       T                     @     �?'             P@       ������������������������       �        !             L@        U       Z                   #@      �?              @        V       Y                    �?      �?             @       W       X                   �>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ]       f                    !@���B�?,           p~@        ^       _                     @r٣����?            �@@        ������������������������       �        	             2@        `       a                    �?��S���?             .@        ������������������������       �                     @        b       c                 03�6@���!pc�?	             &@        ������������������������       �                      @        d       e                    �?�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        g                         @S@8R����?           `|@       h                          @߷���?           P|@       i       l                    ,@������?           �{@        j       k                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        m       �                     �?��#:���?           �{@        n       �                    �?��}*_��?2            @T@       o       �                    �?$��m��?0            �S@       p       q                   �9@�w�r��?/            @S@        ������������������������       �                     &@        r       �                    �?����e��?)            �P@       s       t                    �?��c:�?             G@        ������������������������       �                     ,@        u       �                    �?     ��?             @@       v       �                    K@d��0u��?             >@       w       �                   �G@R�}e�.�?             :@       x       �                 `f�D@�q�q�?             5@       y       �                 �TaA@�d�����?
             3@       z       �                   �E@     ��?	             0@       {       �                   �>@8�Z$���?             *@       |       }                   �;@�8��8��?             (@        ������������������������       �                     @        ~                        03k:@�����H�?             "@        ������������������������       �                      @        �       �                 `fF<@؇���X�?             @       ������������������������       �z�G�z�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                    L@��Q��?             4@       �       �                    �?�����?             3@        �       �                 @�pX@�q�q�?             @       �       �                 ���S@�q�q�?             @        ������������������������       �                     �?        �       �                 ��hU@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �D@�	j*D�?             *@        �       �                    7@�q�q�?             @        ������������������������       �                     �?        �       �                 ���M@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �                          �?�:k �:�?�            pv@       �       �                    @@�)���?�            u@       �       �                    �?��POc�?�            @p@        �       �                   �6@�+$�jP�?             ;@        �       �                    5@      �?             @       �       �                 �{@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   @@���}<S�?             7@       �       �                 ���@r�q��?	             (@        ������������������������       �                     @        �       �                   @<@�<ݚ�?             "@       ������������������������       �����X�?             @        ������������������������       �                      @        ������������������������       �                     &@        �       �                   �>@ �����?�             m@       �       �                 0��D@�#-���?            @j@       �       �                     @�b�E�V�?|            �i@        ������������������������       �                     ?@        �       �                   �<@���	D�?g            �e@       �       �                    �?|E+�	��?_            @d@       �       �                 ���@ 	��p�?S             b@        �       �                 ���@      �?              @       �       �                    �?؇���X�?             @        ������������������������       �                     �?        �       �                    :@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �3@A_�&�?M             a@        �       �                 ��Y @      �?             8@       �       �                    1@d}h���?	             ,@        �       �                 pf�@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �2@"pc�
�?             &@        ������������������������       �                     �?        �       �                 �?�@z�G�z�?             $@       ������������������������       �                     @        ������������������������       �      �?             @        ������������������������       �                     $@        �       �                   �:@ \sF��?=            @\@        ������������������������       �                    �E@        �       �                    �?@4և���?'            �Q@        �       �                 ��(@�IєX�?             1@       �       �                  s�@$�q-�?	             *@        ������������������������       �                      @        ������������������������       ��C��2(�?             &@        ������������������������       �                     @        �       �                   �;@�NW���?            �J@        ������������������������       �                     @        �       �                   @<@p���?             I@       �       �                 ��) @@�E�x�?            �H@       ������������������������       �                    �C@        �       �                 pf� @ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     �?        �       �                   �8@@�0�!��?             1@        �       �                    5@ףp=
�?             $@        �       �                  s�@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �&B@����X�?             @        ������������������������       �                     �?        �       �                    �?r�q��?             @       ������������������������       �                     @        �       �                    ;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�θ�?             *@        ������������������������       �                     �?        �       �                 ���"@r�q��?             (@       ������������������������       �                      @        �       �                 ���)@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                     @      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        �       �                    �?
;&����?             7@       �       �                     @�G��l��?             5@        ������������������������       �                     �?        �       �                 �!B@      �?             4@       �       �                 ��I @�q�q�?
             .@       �       �                    �?�eP*L��?             &@        ������������������������       �                     @        �       �                   �@      �?              @        ������������������������       �                     @        �       �                 �?�@���Q��?             @        ������������������������       �                     �?        �       �                   �?@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @                                 �N@�kb97�?/            @S@                               �E@ �q�q�?+             R@                             `fF)@t��ճC�?             F@             
                @3�@(;L]n�?             >@                                �B@$�q-�?	             *@        ������������������������       �                     @                                 �?؇���X�?             @        ������������������������       �                      @              	                  �C@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             1@                                 �?؇���X�?             ,@        ������������������������       �                     @                              03�2@"pc�
�?             &@                               @D@      �?             @                               @B@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     <@                                  @z�G�z�?             @                                �P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     6@        ������������������������       �                     $@        ������������������������       �                     �?        �t�bh�h*h-K ��h/��R�(KMKK��h]�B�       0|@     Pp@      N@     �d@      @     �E@              A@      @      "@      @      @              @      @       @      @                       @               @      L@     �^@     �G@     �N@     �@@      M@      @     �@@              �?      @      @@      @      ?@               @      @      7@      �?      2@      �?      @      �?      @               @      �?      �?              @              (@      @      @              @      @      �?      @                      �?       @      �?              �?       @              ;@      9@      7@      7@      0@      @              �?      0@      @      .@      @       @              *@      @      @      @               @      @      @      @      �?       @              @      �?       @      �?              �?       @               @                       @      @              �?              @      1@      @      1@      @      *@       @      &@              &@       @              @       @      @                       @              @      �?              @       @      �?       @      �?                       @      @              ,@      @      @              $@      @               @      $@      �?      �?      �?      �?                      �?      "@              "@     �N@      @     �N@              L@      @      @      @      �?      �?      �?      �?                      �?       @                      @      @             px@      X@       @      9@              2@       @      @              @       @      @               @       @      �?       @                      �?     �w@     �Q@     �w@     �Q@     Pw@     �Q@      �?       @      �?                       @     @w@      Q@     �I@      >@     �I@      ;@     �I@      :@      &@              D@      :@      ;@      3@      ,@              *@      3@      &@      3@      @      3@      @      ,@      @      ,@      @      &@       @      &@      �?      &@              @      �?       @               @      �?      @      �?      @               @      �?              @                      @       @                      @      @               @              *@      @      *@      @      @       @      �?       @              �?      �?      �?      �?                      �?      @              "@      @       @      @      �?              �?      @              @      �?              @                      �?              �?              @     t@      C@     �r@      C@     @l@      A@      6@      @      �?      @      �?      �?      �?                      �?               @      5@       @      $@       @      @              @       @      @       @       @              &@             �i@      =@      h@      2@     �g@      0@      ?@             �c@      0@     �b@      *@     �`@      $@      @       @      @      �?      �?              @      �?      @                      �?              �?      `@       @      5@      @      &@      @       @      �?       @                      �?      "@       @      �?               @       @      @               @       @      $@              [@      @     �E@             @P@      @      0@      �?      (@      �?       @              $@      �?      @             �H@      @              @     �H@      �?      H@      �?     �C@              "@      �?              �?      "@              �?              ,@      @      "@      �?       @      �?       @                      �?      @              @       @              �?      @      �?      @              �?      �?      �?                      �?      $@      @              �?      $@       @       @               @       @               @       @               @       @      �?              �?       @      (@      &@      $@      &@              �?      $@      $@      $@      @      @      @      @              @      @              @      @       @      �?               @       @              �?       @      �?      @                      @       @             @R@      @     @Q@      @     �D@      @      =@      �?      (@      �?      @              @      �?       @              @      �?              �?      @              1@              (@       @      @              "@       @       @       @       @      �?      �?      �?      �?                      �?      @              <@              @      �?      �?      �?              �?      �?              @              6@              $@                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ��hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM+huh*h-K ��h/��R�(KM+��h|�B�J         |                  �#@T�����?�           @�@                                   +@X�.;v��?�            �q@        ������������������������       �                     @               I                 ���@�L�w��?�            �q@              H                 0�w@�:���?\             a@              !                 pff@�6���?Z            �`@                                   �?0)RH'�?1            @Q@              	                     @     8�?/             P@        ������������������������       �                     &@        
                          �2@ {��e�?(            �J@        ������������������������       �                      @                                  @<@@�0�!��?&            �I@                                  �?�������?             A@                                   �?      �?
             (@        ������������������������       �                     @                                  �7@      �?              @                                ���@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                  �:@r�q��?             @        ������������������������       �                     �?                                ���@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �      �?             @                                   �?��2(&�?             6@        ������������������������       �                     @                                  �7@�S����?             3@        ������������������������       �                     "@                                ��@�z�G��?             $@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     1@        ������������������������       �                     @        "       #                   �4@�	j*D�?)            @P@        ������������������������       �                     "@        $       -                    �?X�Cc�?#             L@        %       ,                    �?     ��?
             0@       &       +                   @B@d}h���?	             ,@       '       *                 ��@8�Z$���?             *@       (       )                 ���@�8��8��?             (@        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        .       7                    �?R���Q�?             D@        /       4                   �<@�����H�?             2@       0       1                  ��@@4և���?	             ,@        ������������������������       �                     @        2       3                 ��(@ףp=
�?             $@       ������������������������       ������H�?             "@        ������������������������       �                     �?        5       6                   �>@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        8       G                    �?�X����?             6@       9       :                 ��@      �?             4@        ������������������������       �                     @        ;       D                 P�N@�q�q�?	             .@       <       A                   �:@�	j*D�?             *@       =       @                   �6@      �?              @        >       ?                 �1@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        B       C                 �?$@���Q��?             @       ������������������������       �      �?             @        ������������������������       �                     �?        E       F                   �:@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        J       K                 �?�@�9��~�?V            �a@        ������������������������       �                     >@        L       U                 pF @p�̔B��?C            @\@        M       P                    :@��S���?
             .@        N       O                 ���@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        Q       R                    �?���|���?             &@        ������������������������       �                     @        S       T                    �?և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        V       {                   �M@�+�$f��?9            �X@       W       z                 `f#@�^'�ë�?8            @X@       X       w                    �?�Ra����?4             V@       Y       v                    �?���W���?2            �U@       Z       u                   @@@�̨�`<�?1            @U@       [       ^                    �?������?'            �Q@        \       ]                 `�X!@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        _       r                 ���"@(��+�?"            �N@       `       a                   �2@�t����?            �I@        ������������������������       �                     (@        b       q                 ���!@8�Z$���?            �C@       c       d                   �3@"pc�
�?            �@@        ������������������������       �                      @        e       f                   �:@��� ��?             ?@        ������������������������       �                     "@        g       j                 ��) @"pc�
�?             6@       h       i                    ?@      �?             0@       ������������������������       �                     .@        ������������������������       �                     �?        k       l                   �;@      �?             @        ������������������������       �                      @        m       p                    >@      �?             @       n       o                 pf� @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        s       t                   �<@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        
             .@        ������������������������       �                     �?        x       y                 @�!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     �?        }       ~                    �?x>ԛ/��?	           �z@        ������������������������       �                     1@               *                   @��3���?           �y@       �       �                   �1@���`��?�             y@        �       �                    @^��>�b�?'            @P@       �       �                    �?,���i�?            �D@       �       �                 P��%@�KM�]�?             C@        ������������������������       �                     �?        �       �                    �?�L���?            �B@       ������������������������       �                     5@        �       �                 ���2@     ��?
             0@       ������������������������       �                     "@        �       �                   �0@և���X�?             @       �       �                 `�I@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   XB@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �? �q�q�?             8@        ������������������������       �                     @        �       �                    �?�IєX�?             1@        ������������������������       �                     @        �       �                    �?�C��2(�?             &@       �       �                    @r�q��?             @        ������������������������       �                      @        �       �                 ��T?@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �                       ���S@Z�cI��?�            u@       �       �                 0#�9@B�Y�9d�?�            �q@        �       �                 ��Y7@OX���?Y            �a@       �       �                    @�X���?R            �`@       �       �                   @I@     ��?P             `@       �       �                 ��6@L
�q��?K            �]@       �       �                 pF%@�����?H            �\@        �       �                 �yW$@�eP*L��?             &@        ������������������������       �                     �?        �       �                   �7@      �?             $@        ������������������������       �                      @        �       �                    @@      �?              @        ������������������������       �                     @        �       �                   @E@      �?             @       �       �                   @A@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�V	�?l�?A            �Y@        �       �                   �:@�G�z�?             D@        �       �                 P�>,@�θ�?             *@       �       �                 ��*@�q�q�?             "@       �       �                     @      �?              @       ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                     @�����H�?             ;@        ������������������������       �                     $@        �       �                   �D@@�0�!��?             1@       �       �                    �?      �?             0@        ������������������������       �                     @        �       �                    �?"pc�
�?	             &@       �       �                    �?z�G�z�?             $@       �       �                 03�1@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �=@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   @<@���N8�?(            �O@       �       �                     @�8��8��?             B@        �       �                   �(@z�G�z�?
             .@        ������������������������       �                     @        �       �                   �9@      �?             (@       ������������������������       �                     @        �       �                    �?���Q��?             @        ������������������������       �                     �?        �       �                   �*@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     5@        ������������������������       �                     ;@        ������������������������       �                     @        �       �                 `f'@ףp=
�?             $@        �       �                   �P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     &@        �       �                    �?������?]            @a@        �       �                     @�����?             E@       ������������������������       �                     C@        ������������������������       �                     @        �                         �J@r�qG�?A             X@       �       �                 `f�:@�^�����?8            �U@        �       �                     �?���Q��?
             .@       �       �                   @G@�<ݚ�?             "@       �       �                   @B@      �?             @        ������������������������       �      �?              @        ������������������������       �      �?              @        ������������������������       �                     @        �       �                    :@�q�q�?             @       �       �                    �?      �?             @        ������������������������       �                     �?        �       �                   �@@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �                         �G@v���EO�?.            �Q@       �                          �?�'�`d�?+            �P@       �                          A@p9W��S�?             C@       �       �                    �?����"�?             =@        �       �                    ?@      �?             @       �       �                 @�J@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �                         �?@�LQ�1	�?             7@       �       �                   �?@����X�?             5@        ������������������������       �                     @        �                       ��?P@r�q��?             2@       �                         �=@d}h���?
             ,@       �                           @�θ�?	             *@       �                           �?�����H�?             "@       �                       ��yC@      �?              @        �                          �A@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@        	                         �? �Cc}�?             <@        
                          �?�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @                              `�iJ@�KM�]�?             3@                               x#J@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     &@                              p"�S@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        	             $@                                 �?����X�?!             L@                               �:@г�wY;�?             A@                                 �?�����H�?             "@        ������������������������       �                     @                              ���i@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     9@                                 �?�X����?             6@        ������������������������       �                      @               !                Ј�U@      �?	             ,@        ������������������������       �                     @        "      )                   �?���|���?             &@       #      (                p"�X@X�<ݚ�?             "@       $      %                   �?r�q��?             @        ������������������������       �                     @        &      '                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �t�b��     h�h*h-K ��h/��R�(KM+KK��h]�B�       0|@     Pp@     `l@      M@              @     `l@     �J@     �Y@      A@     �Y@      ?@      M@      &@     �J@      &@      &@              E@      &@               @      E@      "@      9@      "@      @      @              @      @       @      �?      �?              �?      �?              @      �?      �?              @      �?      �?              @      �?      3@      @      @              0@      @      "@              @      @              @      @              1@              @             �F@      4@      "@              B@      4@      @      &@      @      &@       @      &@      �?      &@              @      �?      @      �?              �?               @              ?@      "@      0@       @      *@      �?      @              "@      �?       @      �?      �?              @      �?              �?      @              .@      @      .@      @      @              $@      @      "@      @      @      �?       @      �?              �?       @              @               @      @       @       @              �?      �?      �?      �?                      �?               @              @      _@      3@      >@             �W@      3@      @       @      @      �?      @                      �?      @      @              @      @      @              @      @             �U@      &@     �U@      $@     �S@      $@     @S@      "@      S@      "@     �N@      "@       @      �?       @                      �?     �J@       @     �F@      @      (@             �@@      @      ;@      @               @      ;@      @      "@              2@      @      .@      �?      .@                      �?      @      @               @      @      �?      �?      �?              �?      �?               @              @               @       @       @                       @      .@              �?              �?      �?      �?                      �?      "@                      �?      l@     `i@              1@      l@     @g@      k@     @g@      <@     �B@      @      B@      @      A@      �?              @      A@              5@      @      *@              "@      @      @      @      �?      @                      �?              @      �?       @      �?                       @      7@      �?      @              0@      �?      @              $@      �?      @      �?       @              @      �?      @                      �?      @             �g@     �b@     �e@     @[@     �X@     �F@     �U@     �F@     �U@     �D@     �S@      D@     �S@      B@      @      @              �?      @      @               @      @      @      @              �?      @      �?      �?              �?      �?                       @     @R@      >@      *@      ;@      $@      @      @      @      @       @      @       @       @                      �?      @              @      8@              $@      @      ,@       @      ,@              @       @      "@       @       @      �?      @              @      �?              �?      @      �?                      @              �?      �?              N@      @     �@@      @      (@      @      @              "@      @      @               @      @      �?              �?      @              @      �?              5@              ;@                      @      "@      �?      �?      �?              �?      �?               @                      @      &@             �R@      P@      @      C@              C@      @             �Q@      :@      N@      :@      @      "@       @      @       @       @      �?      �?      �?      �?              @      @       @       @       @      �?              �?       @               @      �?               @              K@      1@      J@      ,@      ;@      &@      2@      &@      @      @      @      �?      @                      �?               @      .@       @      .@      @              @      .@      @      &@      @      $@      @       @      �?      @      �?      �?      �?      �?                      �?      @              �?               @       @      �?              @                       @      "@              9@      @       @      �?              �?       @              1@       @      @       @      @                       @      &@               @      @              @       @              $@              0@      D@      �?     �@@      �?       @              @      �?      @      �?                      @              9@      .@      @       @              @      @      @              @      @      @      @      �?      @              @      �?      �?              �?      �?              @                       @       @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ��nhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM!huh*h-K ��h/��R�(KM!��h|�B@H                            @�"Y�\7�?�           @�@              Y                    �?��d1h��?�           �@               X                    @��Hg���?�             l@              G                   �>@�GN�z�?�            �k@              @                    @&���7��?c            `b@                                  �?V�L��?\            �`@                                    @     ��?             @@        ������������������������       �        
             1@        	       
                   �+@�q�q�?
             .@        ������������������������       �                     @                                   �?X�<ݚ�?             "@                                  :@և���X�?             @        ������������������������       �                      @                                   �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @               !                     @�t����?H            �Y@                                   �?ףp=
�?              D@                                  2@Pa�	�?            �@@                                ��Y)@؇���X�?             @        ������������������������       �                     @                                   :@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     :@                                   �?և���X�?             @        ������������������������       �                     �?                                     �?      �?             @                               ���`@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        "       ?                    �?�P�*�?(             O@       #       :                    �?Ɣ��Hr�?%            �M@       $       5                   �9@�L�lRT�?            �F@       %       &                 ��}@�5��?             ;@        ������������������������       �                     @        '       ,                    3@�q�q�?             8@        (       +                    $@�8��8��?             (@        )       *                   �&@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        -       4                 pff@�q�q�?	             (@       .       /                 ���@����X�?             @        ������������������������       �                     @        0       1                    �?      �?             @        ������������������������       �                     �?        2       3                   �7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        6       7                 @3�@�E��ӭ�?             2@       ������������������������       �                     $@        8       9                 @3#%@      �?              @       ������������������������       �                     @        ������������������������       �                     @        ;       <                 `f�-@      �?
             ,@        ������������������������       �                     @        =       >                 @3�/@�z�G��?             $@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        A       B                 ��	5@8�Z$���?             *@        ������������������������       �                     �?        C       D                   �0@�8��8��?             (@       ������������������������       �                     $@        E       F                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        H       I                 ��n @F��}��?.            @R@        ������������������������       �                     �?        J       W                    �? �q�q�?-             R@       K       L                    �?��<D�m�?            �H@       ������������������������       �                     ;@        M       N                    �?��2(&�?             6@        ������������������������       �                     @        O       P                 ��Y.@z�G�z�?
             .@        ������������������������       �                      @        Q       V                     @$�q-�?             *@       R       U                    6@ףp=
�?             $@        S       T                   �@@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     7@        ������������������������       �                     @        Z       ]                    @�\���?           |@        [       \                     @�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ^       �                  x#J@�7�WR�?           �{@       _       �                     �?�+�$f��?�            �x@        `       �                    �?�����?#            �H@       a       b                   �;@�q�q�?"             H@        ������������������������       �                     �?        c       �                    �?��k=.��?!            �G@       d                           R@z�G�z�?            �F@       e       ~                   �L@"pc�
�?             F@       f       k                   @=@x�����?            �C@        g       h                   �G@��S�ۿ?	             .@       ������������������������       �                     &@        i       j                    J@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        l       q                    �?�q�q�?             8@        m       n                    A@�q�q�?             @        ������������������������       �                     �?        o       p                    G@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        r       y                   �<@���N8�?             5@       s       t                   �>@�	j*D�?             *@        ������������������������       �                      @        u       v                   �A@"pc�
�?             &@        ������������������������       �                     @        w       x                 ��yC@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        z       {                   �H@      �?              @       ������������������������       �                     @        |       }                   �J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                     @�4rU��?�            pu@        �       �                    :@ ���g=�?.            @Q@       �       �                   @A@�r����?'             N@       �       �                    �?tk~X��?             B@       �       �                    @@r�q��?             >@       �       �                 `��,@ȵHPS!�?             :@       �       �                    �?؇���X�?             5@        ������������������������       �                     �?        �       �                    &@ףp=
�?             4@       �       �                   �6@r�q��?             (@        ������������������������       ��q�q�?             @        ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �      �?             @        �       �                   �7@�q�q�?             @        ������������������������       �                     @        �       �                   �<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 `f'@ �q�q�?             8@        �       �                   @H@z�G�z�?             @        ������������������������       �                     @        �       �                   �P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     3@        ������������������������       �                     "@        �       �                 ��y @���	���?�             q@       �       �                    �?Xny��?u            �f@        �       �                 ���@$�q-�?            �C@        �       �                    9@�����H�?             2@        �       �                    �?      �?             @       �       �                 ��y@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        
             ,@        �       �                   �=@���N8�?             5@       �       �                  ��@��S�ۿ?
             .@        ������������������������       �                      @        �       �                 ��(@$�q-�?             *@       �       �                    �?�8��8��?             (@       ������������������������       ��C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ��) @      �?Y             b@       �       �                 �?�@�Z��L��?X            �a@       �       �                 ���@ 	��p�?5            �U@        �       �                 ���@�S����?             3@       �       �                    �?�����H�?             2@       �       �                   �>@؇���X�?
             ,@        �       �                    :@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                 �{@ =[y��?)             Q@       �       �                 ���@��p\�?            �D@       ������������������������       �                     :@        �       �                 P�N@z�G�z�?             .@       �       �                 �?$@r�q��?             (@       �       �                    ;@z�G�z�?             $@        ������������������������       �                     @        �       �                   �=@����X�?             @        ������������������������       ����Q��?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    :@�q�q�?             @        ������������������������       �                     �?        �       �                    D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ;@        �       �                    �?"pc�
�?#            �K@       �       �                 @3�@�����?!            �H@        �       �                    �?և���X�?             @       �       �                   �?@      �?             @        ������������������������       �                     �?        �       �                   �D@���Q��?             @       �       �                   �A@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �1@؇���X�?             E@        ������������������������       ��q�q�?             @        �       �                   �3@��-�=��?            �C@        ������������������������       �����X�?             @        �       �                    ?@      �?             @@       ������������������������       �                     7@        �       �                   �@@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                    ,@0�>���?3            �V@        �       �                 �y.@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �? p�/��?1            @V@       �       �                    �? Df@��?,            �T@       �       �                    �?�g�y��?#             O@        �       �                 `v�0@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �<@P����?!            �M@       ������������������������       �                    �D@        �       �                 ���"@�X�<ݺ?             2@       ������������������������       �                     $@        �       �                 ��Y)@      �?              @        �       �                    ?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             5@        �       �                    �?�q�q�?             @        �       �                  �v6@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �                          �?     ��?             H@       �                          �5@������?             >@        ������������������������       �                      @                              `f�N@d}h���?             <@        ������������������������       �                     ,@              
                    �?և���X�?             ,@                             03�U@�q�q�?             (@        ������������������������       �                     @              	                   �?�����H�?             "@                              p�w@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @                                 �?�E��ӭ�?             2@                                 6@���Q��?             @        ������������������������       �                      @                                 �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                 �?8�Z$���?	             *@        ������������������������       �                     @                                @F@      �?              @                                �;@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @                                  @�}�+r��?             C@                                �?�C��2(�?             6@                              ���3@      �?              @        ������������������������       �                     �?                              ��T?@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     ,@        ������������������������       �        	             0@        �t�bh�h*h-K ��h/��R�(KM!KK��h]�B       �|@     `o@     �z@      o@     �K@     @e@      I@     @e@      G@     @Y@     �A@     �X@      @      ;@              1@      @      $@              @      @      @      @      @               @      @       @               @      @               @              >@      R@      @      B@      �?      @@      �?      @              @      �?      @      �?                      @              :@      @      @              �?      @      @      @      �?              �?      @                       @      :@      B@      7@      B@      0@      =@      &@      0@      @               @      0@      �?      &@      �?       @      �?                       @              "@      @      @       @      @              @       @       @      �?              �?       @               @      �?              @              @      *@              $@      @      @      @                      @      @      @      @              @      @              @      @              @              &@       @              �?      &@      �?      $@              �?      �?      �?                      �?      @     @Q@      �?              @     @Q@      @      G@              ;@      @      3@              @      @      (@       @              �?      (@      �?      "@      �?       @      �?                       @              @              @              7@      @              w@     �S@      �?       @               @      �?             w@     �Q@     �u@      F@     �C@      $@      C@      $@              �?      C@      "@      B@      "@      B@       @      ?@       @      ,@      �?      &@              @      �?              �?      @              1@      @      �?       @              �?      �?      �?      �?                      �?      0@      @      "@      @               @      "@       @      @              @       @               @      @              @      �?      @              �?      �?              �?      �?              @                      �?       @              �?             Ps@      A@     �N@       @      J@       @      =@      @      9@      @      7@      @      2@      @              �?      2@       @      $@       @      �?       @      "@               @              @               @       @      @       @      @              �?       @      �?                       @      7@      �?      @      �?      @              �?      �?              �?      �?              3@              "@              o@      :@     @d@      5@      B@      @      0@       @       @       @      �?       @      �?                       @      �?              ,@              4@      �?      ,@      �?       @              (@      �?      &@      �?      $@      �?      �?              �?              @             �_@      2@     �_@      0@     @T@      @      0@      @      0@       @      (@       @      @       @      @                       @       @              @                      �?     @P@      @      C@      @      :@              (@      @      $@       @       @       @      @              @       @      @       @       @               @               @      �?      �?              �?      �?              �?      �?              ;@             �F@      $@     �C@      $@      @      @      @      @              �?      @       @      @      �?       @      �?      �?                      �?              �?      B@      @      �?       @     �A@      @      @       @      >@       @      7@              @       @               @      @              @                       @     �U@      @      �?      �?              �?      �?             @U@      @     @T@       @      N@       @       @      �?       @                      �?      M@      �?     �D@              1@      �?      $@              @      �?      �?      �?              �?      �?              @              5@              @       @      �?       @      �?                       @      @              5@      ;@       @      6@       @              @      6@              ,@      @       @      @       @      @              �?       @      �?       @      �?                       @              @       @              *@      @       @      @               @       @      �?              �?       @              &@       @      @              @       @       @       @       @                       @      @              B@       @      4@       @      @       @              �?      @      �?      @                      �?      ,@              0@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJXk�hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM?huh*h-K ��h/��R�(KM?��h|�B�O         �                     @��ے@R�?�           @�@                                   /@�r�����?�            Ps@               
                     �?�C��2(�?             6@                                   �?�<ݚ�?             "@        ������������������������       �                     �?               	                    �?      �?              @                                ���`@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        
             *@               Q                     �?�!I���?�            �q@              P                    @���;+"�?`            �c@              +                   �?@"+q��?_            @c@                                  �;@     ��?&             P@                                   2@      �?             4@        ������������������������       �                     @                                   �?�t����?             1@                                  �?$�q-�?
             *@                                 �6@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @                                   �?���|���?             F@        ������������������������       �                     @                                   �?���"͏�?            �B@        ������������������������       �                      @               *                   @K@8^s]e�?             =@              )                    �?������?             ;@              (                 ��yC@8����?             7@               !                 `fF:@     ��?	             0@        ������������������������       �                     @        "       '                   �A@�q�q�?             (@       #       &                   �>@      �?             $@       $       %                 `f�<@����X�?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ,       3                    �?$�ݏ^��?9            �V@        -       2                    �?@�E�x�?            �H@       .       1                 �D�E@`2U0*��?             9@        /       0                    �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     2@        ������������������������       �                     8@        4       O                  D�\@�4F����?            �D@       5       6                   �9@�d�����?             C@        ������������������������       �                     @        7       >                    D@:ɨ��?            �@@        8       9                    �?؇���X�?             @        ������������������������       �                     �?        :       ;                    �?r�q��?             @        ������������������������       �                     @        <       =                   @B@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ?       H                    �?8�Z$���?             :@        @       G                   �J@      �?              @       A       B                    �?r�q��?             @        ������������������������       �                      @        C       F                    �?      �?             @       D       E                   �H@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        I       N                    �?�X�<ݺ?             2@       J       M                   �J@�C��2(�?             &@        K       L                   �H@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        R       �                    �?��>^�?Q             `@       S       �                   �I@���U��?9            @W@       T       Y                    �?l�Ӑ���?4            �U@        U       V                    4@      �?              @        ������������������������       �                     �?        W       X                 pf�,@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        Z       }                   @D@�2��?0            �S@       [       ^                   �7@.��<�?*            �P@        \       ]                    �?@4և���?	             ,@       ������������������������       �                     *@        ������������������������       �                     �?        _       z                    �?�q����?!            �J@       `       w                    �?�t����?            �I@       a       v                   @A@8����?             G@       b       q                   �@@�99lMt�?            �C@       c       h                    �?�t����?             A@        d       e                   �'@"pc�
�?             &@        ������������������������       �                      @        f       g                    :@�<ݚ�?             "@        ������������������������       �      �?             @        ������������������������       �                     @        i       j                 `fF)@�nkK�?             7@       ������������������������       �                     *@        k       p                   �3@ףp=
�?             $@       l       m                   �;@�����H�?             "@        ������������������������       �                     @        n       o                    =@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        r       s                   �'@z�G�z�?             @        ������������������������       �                      @        t       u                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        x       y                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        {       |                   `A@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ~                          �F@�q�q�?             (@        ������������������������       �                     @        �       �                    �?����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?      �?             B@        �       �                    �?�X�<ݺ?             2@       �       �                   �;@�����H�?             "@        �       �                 ��m1@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        �       �                    �?�X�<ݺ?             2@       �       �                    �?��S�ۿ?             .@       �       �                    �?�C��2(�?	             &@        ������������������������       �                     @        �       �                   �<@؇���X�?             @        ������������������������       �                     @        �       �                   �7@      �?             @        ������������������������       �                     �?        �       �                   �B@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?h�*���?           0y@        �       �                   �7@�Jl$G��?D            �[@        �       �                    @��>4և�?             <@        ������������������������       �                     @        �       �                 �n6@r�q��?             8@       �       �                    �?��Q��?             4@       �       �                 03�@ҳ�wY;�?
             1@        ������������������������       �                      @        �       �                    �?������?             .@       �       �                    �?���|���?             &@       �       �                   �2@�<ݚ�?             "@       ������������������������       �                     @        �       �                   �5@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                 ��&@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                 �?�-@ؤ�u��?3            �T@       �       �                    >@ٜSu��?(            @Q@       �       �                    �?�ɞ`s�?#            �N@       �       �                   �:@�q�q�?!            �L@        ������������������������       �                     @        �       �                    �?H(���o�?            �J@        �       �                    �?�+e�X�?             9@        ������������������������       �                     @        �       �                 ���@�����?             5@        ������������������������       �                     @        �       �                   �<@؇���X�?	             ,@       �       �                   @@$�q-�?             *@       �       �                   @<@r�q��?             @       ������������������������       �z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?���>4��?             <@        ������������������������       �                     (@        �       �                  s�@      �?	             0@        ������������������������       �                     @        �       �                 ��(@�C��2(�?             &@       ������������������������       ������H�?             "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                 03�7@և���X�?             ,@       �       �                    �?�q�q�?	             (@       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                    @����s�?�            @r@        �       �                     @D�n�3�?             3@        �       �                    �?X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @        �       �                 ��T?@�z�G��?             $@        ������������������������       �                     @        �       �                    �?���Q��?             @        ������������������������       �                      @        �       �                     @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       0                  @B@��yP��?�            q@       �       /                   @��^���?�             m@       �       &                   �?.P�'z�?�            `k@       �       �                    �?��SK�?}            �g@        �       �                   �>@      �?             D@       �       �                    �?">�֕�?            �A@       �       �                 ���@$��m��?             :@        ������������������������       �                     @        �       �                    ;@�GN�z�?             6@       �       �                   �9@�	j*D�?             *@       �       �                 @�"@"pc�
�?	             &@       �       �                    5@�����H�?             "@        ������������������������       �                     @        �       �                 pff@z�G�z�?             @        �       �                   �7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    4@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                 @3#%@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        �       �                 ���)@�<ݚ�?             "@        ������������������������       �                     @        �       �                    ;@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                 03�1@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �                         �8@*~k���?a            �b@        �       �                 @3�@ pƵHP�?#             J@       ������������������������       �                     @@        �                          �?P���Q�?             4@       �                         �0@�}�+r��?             3@        �                        �̌!@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     0@        ������������������������       �                     �?                                �;@fhK�4�?>            �X@                              ��@      �?
             0@        ������������������������       �                     @                                 �?�q�q�?             (@                             �@@�<ݚ�?             "@       	      
                  �:@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?                                 �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?              %                   �?��Lɿ��?4            �T@             "                �T�C@ȵHPS!�?0            �S@                              sW@���;QU�?-            @R@                              P��@؇���X�?	             5@       ������������������������       �                     "@                                �=@      �?             (@        ������������������������       �      �?             @        ������������������������       �                     @                              �?�@ ��WV�?$             J@        ������������������������       �                     7@              !                  �?@ 	��p�?             =@                                 >@�����?             5@                             ��) @P���Q�?             4@        ������������������������       �                     &@                              pf� @�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        #      $                   >@z�G�z�?             @       ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        '      .                   �?����X�?             <@       (      -                ���5@���Q��?             4@        )      *                  �*@�����H�?             "@        ������������������������       �                     @        +      ,                  �=@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                      @        ������������������������       �                     *@        1      >                   �?������?            �D@       2      7                   �?�IєX�?             A@        3      6                   @z�G�z�?             @       4      5                   I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        8      9                  �E@XB���?             =@        ������������������������       �        	             .@        :      ;                P�@@4և���?
             ,@        ������������������������       �                     @        <      =                  �F@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �t�bh�h*h-K ��h/��R�(KM?KK��h]�B�       �|@     �o@     �b@     �c@       @      4@       @      @              �?       @      @       @       @               @       @                      @              *@     �b@     @a@     �P@      W@      O@      W@     �@@      ?@      @      .@              @      @      (@      �?      (@      �?       @      �?                       @              @      @              <@      0@              @      <@      "@       @              4@      "@      4@      @      0@      @      "@      @      @              @      @      @      @       @      @       @      @              �?      @                       @      @              @                       @      =@     �N@      �?      H@      �?      8@      �?      @      �?                      @              2@              8@      <@      *@      <@      $@      @              7@      $@      �?      @              �?      �?      @              @      �?       @      �?                       @      6@      @      @      @      @      �?       @              @      �?       @      �?              �?       @              �?                       @      1@      �?      $@      �?       @      �?       @                      �?       @              @                      @      @             �T@      G@     @P@      <@     �M@      <@      @      @              �?      @      @              @      @             �K@      8@      I@      1@      *@      �?      *@                      �?     �B@      0@      B@      .@      @@      ,@      9@      ,@      8@      $@       @      "@               @       @      @       @       @              @      6@      �?      *@              "@      �?       @      �?      @              @      �?              �?      @              �?              �?      @               @      �?       @               @      �?              @              @      �?              �?      @              �?      �?              �?      �?              @      @              @      @       @               @      @              @              2@      2@      �?      1@      �?       @      �?      @              @      �?                      @              "@      1@      �?      ,@      �?      $@      �?      @              @      �?      @              @      �?      �?               @      �?              �?       @              @              @             @s@     �W@     �P@      F@      &@      1@              @      &@      *@      @      *@      @      &@       @              @      &@      @      @       @      @              @       @      @       @                      @       @                      @      �?       @      �?                       @      @              L@      ;@      I@      3@      E@      3@      C@      3@      @              A@      3@      3@      @              @      3@       @      @              (@       @      (@      �?      @      �?      @      �?      �?              @                      �?      .@      *@              (@      .@      �?      @              $@      �?       @      �?       @              @               @              @       @      @       @               @      @               @              n@     �I@      &@       @      @      @      @                      @      @      @      @               @      @               @       @      �?       @                      �?     �l@     �E@     �g@     �D@     @f@     �D@     �c@     �@@      9@      .@      8@      &@      1@      "@              @      1@      @      "@      @      "@       @       @      �?      @              @      �?       @      �?              �?       @               @              �?      �?              �?      �?                       @       @      �?       @                      �?      @       @      @               @       @       @                       @      �?      @              @      �?             �`@      2@     �I@      �?      @@              3@      �?      2@      �?       @      �?      �?      �?      �?              0@              �?             �T@      1@       @       @              @       @      @      @       @      @      �?      @                      �?              �?      �?       @               @      �?             �R@      "@     @Q@      "@      Q@      @      2@      @      "@              "@      @      @      @      @              I@       @      7@              ;@       @      3@       @      3@      �?      &@               @      �?              �?       @                      �?       @              �?      @      �?       @               @      @              4@       @      (@       @      �?       @              @      �?      @      �?                      @      &@               @              *@             �C@       @      @@       @      @      �?      �?      �?      �?                      �?      @              <@      �?      .@              *@      �?      @              @      �?              �?      @              @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ0��JhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM-huh*h-K ��h/��R�(KM-��h|�B@K         x                     @�d��Pb�?�           @�@                                   /@~����m�?�            u@        ������������������������       �                     5@                                   �?�j����?�            �s@                                    �?����}��?K            �_@       ������������������������       �        +             R@                                   �? �Jj�G�?             �K@       ������������������������       �                     @@        	                           6@�nkK�?             7@        
                           �?�C��2(�?             &@        ������������������������       �                     @                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             (@               5                 ��D:@�3�B���?v            �g@               4                    M@$��$�L�?5            �S@              #                   �<@�:�^���?4            �S@               "                    �?�ݜ�?            �C@                                  @$G$n��?            �B@        ������������������������       �                      @                                  �'@д>��C�?             =@                                  �1@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               !                 `��,@PN��T'�?             ;@                                 �;@��s����?             5@       ������������������������       �                     0@                                  �*@z�G�z�?             @        ������������������������       �                     @                                 ��\+@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        $       3                   @E@�7��?            �C@       %       &                     �? 	��p�?             =@        ������������������������       �                     @        '       2                   @D@HP�s��?             9@       (       )                   �@@���N8�?             5@        ������������������������       �                      @        *       1                    �?$�q-�?	             *@       +       ,                   �'@ףp=
�?             $@        ������������������������       �                     @        -       0                   �3@r�q��?             @       .       /                   @B@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �      �?             @        ������������������������       �                     $@        ������������������������       �                     �?        6       k                    �?��N`.�?A            �[@       7       L                    �?���ȫ�?4            �T@        8       K                     �?�n_Y�K�?             :@       9       F                 �D�G@�q�q�?             8@       :       A                    ?@��
ц��?             *@        ;       @                    =@z�G�z�?             @       <       ?                 03SA@      �?             @       =       >                 �ܵ<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        B       E                   �L@      �?              @       C       D                   �B@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        G       H                 @�pX@�C��2(�?             &@       ������������������������       �                     "@        I       J                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        M       b                    �?���X�?$             L@       N       _                   @J@�����?             C@       O       X                   �?@�5��?             ;@       P       W                     �?������?             1@       Q       V                   �>@������?
             .@        R       S                   �;@z�G�z�?             @        ������������������������       �                     �?        T       U                 `fF<@      �?             @        ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �                      @        Y       ^                 `f?@�z�G��?             $@       Z       [                   �E@      �?              @        ������������������������       �                     @        \       ]                   @G@z�G�z�?             @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                      @        `       a                    R@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        c       h                   �G@r�q��?             2@       d       g                    =@��S�ۿ?
             .@        e       f                   �9@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        i       j                 ���W@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        l       w                     �?�>4և��?             <@       m       v                   �B@��<b���?             7@       n       u                   �d@�n_Y�K�?             *@       o       r                   �<@      �?              @        p       q                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        s       t                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                     @        y       �                    �?b����o�?�            pw@        z       �                    �?��e�B��?E            �Y@       {       �                    �?L�qA��?3            �R@        |       �                    �?�q�q�?             8@        }       ~                   �+@      �?              @        ������������������������       �                     @               �                   �6@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                 Ь* @     ��?             0@       �       �                    4@"pc�
�?	             &@        �       �                    1@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                    9@      �?              @        ������������������������       �                     �?        �       �                 ���@؇���X�?             @        ������������������������       �                     @        ������������������������       ��q�q�?             @        �       �                 03�'@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?j���� �?             �I@       �       �                    @     ��?             @@       �       �                   @B@��>4և�?             <@       �       �                    �?�q�q�?             8@       �       �                    0@8����?             7@        ������������������������       �                     �?        �       �                    �?���!pc�?             6@       �       �                   �@������?             1@       �       �                 ���@$�q-�?             *@       ������������������������       �                     @        �       �                 �&B@r�q��?             @       �       �                    4@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                 ��&@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �:@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   #@      �?             @        ������������������������       �                     �?        �       �                    �?�q�q�?             @       �       �                    I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                     @�\��N��?             3@       �       �                   �>@     ��?	             0@       �       �                    �?�q�q�?             (@        �       �                    -@      �?             @       �       �                   �&@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                    -@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �<@�q�q�?             ;@       �       �                    �?�û��|�?             7@        �       �                    �?�q�q�?             (@        �       �                 `�@1@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    :@և���X�?             @       �       �                    @z�G�z�?             @        ������������������������       �                      @        �       �                    1@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                 ���3@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     @        �                          �?Dg�-N�?�            q@       �                          �?4��?�?�             j@       �       �                    �?@��Y��?�            �i@        �       �                    ;@���.�6�?             G@        �       �                 0S�*@����X�?             @       �       �                   �4@r�q��?             @       �       �                   �3@�q�q�?             @        ������������������������       �                     �?        �       �                 �{@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                 ���@ ���J��?            �C@        �       �                 ���@      �?
             0@       ������������������������       �                     (@        �       �                    =@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     7@        �                       �T)D@$��$�L�?e            �c@       �                         @@@�:�]��?a             c@       �                         �?@L�'�7��?I            @]@       �       �                 @33@�L���?E            �[@        �       �                    6@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 @3�@��Wv��?C             [@        �       �                 �?$@@3����?             K@        �       �                   �:@���7�?             6@       ������������������������       �                     ,@        �       �                 ��@      �?              @        ������������������������       �                      @        �       �                   �=@r�q��?             @       ������������������������       �      �?             @        ������������������������       �                      @        ������������������������       �                     @@        �       �                 ���!@�����H�?$             K@       �       �                 ��) @     ��?             @@       �       �                    4@HP�s��?             9@        �       �                   �1@���Q��?             @        ������������������������       ��q�q�?             @        ������������������������       �      �?              @        ������������������������       �                     4@        �       �                 pf� @և���X�?             @        ������������������������       �                     �?        �       �                   �7@�q�q�?             @        ������������������������       �                     @        �       �                   �;@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 ���"@���7�?             6@        ������������������������       �                      @                               ���#@@4և���?             ,@                               �<@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @                              P�@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @              	                  �E@������?             B@       ������������������������       �                     6@        
                      @3�@@4և���?
             ,@                             ��Y@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @                                 >@z�G�z�?             @        ������������������������       ��q�q�?             @        ������������������������       �                      @                              ���*@      �?             @        ������������������������       �                     �?        ������������������������       �                     @                                 �?��ɉ�?*            @P@                                 �?h�����?             <@                                 �?r�q��?             @        ������������������������       �                     @                               �v6@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     6@              ,                   $@���@��?            �B@              #                   @���Q��?             4@                                  �?      �?              @        ������������������������       �                     @        !      "                   @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        $      '                   @�q�q�?             (@       %      &                   �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        (      )                   �?�q�q�?             @        ������������������������       �                     @        *      +                03�;@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     1@        �t�b�     h�h*h-K ��h/��R�(KM-KK��h]�B�       @{@     @q@     @b@     �g@              5@     @b@     @e@      �?     �_@              R@      �?      K@              @@      �?      6@      �?      $@              @      �?      @      �?                      @              (@      b@      F@     �Q@       @     �Q@      @      A@      @      @@      @       @              8@      @      �?      �?      �?                      �?      7@      @      1@      @      0@              �?      @              @      �?      �?      �?                      �?      @               @             �B@       @      ;@       @      @              7@       @      4@      �?       @              (@      �?      "@      �?      @              @      �?       @      �?      �?      �?      �?              @              @              @      �?      $@                      �?     �R@      B@     �I@      ?@      $@      0@       @      0@      @      @      @      �?      @      �?      �?      �?      �?                      �?       @              �?              @      @       @      @              @       @              �?              �?      $@              "@      �?      �?              �?      �?               @             �D@      .@      :@      (@      0@      &@      *@      @      &@      @      �?      @              �?      �?      @      �?      �?               @      $@               @              @      @      �?      @              @      �?      @      �?      �?              @       @              $@      �?      $@                      �?      .@      @      ,@      �?      @      �?      @                      �?      &@              �?       @      �?                       @      7@      @      2@      @       @      @      @      @       @      �?       @                      �?      �?      @      �?                      @      @              $@              @              r@     @U@      G@      L@      <@     �G@      @      1@       @      @              @       @       @       @                       @      @      &@       @      "@      �?       @               @      �?              �?      @              �?      �?      @              @      �?       @      @       @      @                       @      5@      >@      &@      5@      &@      1@       @      0@      @      0@      �?              @      0@      @      *@      �?      (@              @      �?      @      �?      @      �?                      @              �?      @      �?      @                      �?       @      @       @                      @      �?              @      �?      �?               @      �?      �?      �?      �?                      �?      �?                      @      $@      "@      @      "@      @      @      �?      @      �?       @      �?                       @              �?      @       @               @      @                      @      @              2@      "@      ,@      "@      @       @      �?      @      �?                      @      @      @      �?      @               @      �?       @      �?                       @       @              $@      �?              �?      $@              @             �n@      =@     �g@      4@      g@      3@     �E@      @      @       @      @      �?       @      �?      �?              �?      �?      �?                      �?      @                      �?      C@      �?      .@      �?      (@              @      �?       @      �?      �?              7@             �a@      0@     �a@      (@     �Z@      &@     �Y@      "@      �?       @      �?                       @     @Y@      @     �J@      �?      5@      �?      ,@              @      �?       @              @      �?      @      �?       @              @@              H@      @      ;@      @      7@       @      @       @       @      �?      �?      �?      4@              @      @              �?      @       @      @              �?       @               @      �?              5@      �?       @              *@      �?      @      �?      @                      �?      @              @       @               @      @             �A@      �?      6@              *@      �?      @      �?      @                      �?      @              �?      @      �?       @               @      @      �?              �?      @              L@      "@      ;@      �?      @      �?      @               @      �?       @                      �?      6@              =@       @      (@       @      @      �?      @              �?      �?              �?      �?              @      @      �?      @      �?                      @      @       @      @              �?       @               @      �?              1@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJڡWhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM1huh*h-K ��h/��R�(KM1��h|�B@L         �                     @�1�uџ�?�           @�@               _                    �?2������?�            �s@              
                    �?և���X�?�            �m@                                  �H@�k~X��?,             R@       ������������������������       �        &             O@               	                    �?ףp=
�?             $@                                   K@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @               *                   �?@Z�J�p�?g            �d@                                    �?�?�'�@�?3             S@                                  �;@�חF�P�?             ?@                                   �?�q�q�?             @                                 �7@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?                                   �?H%u��?             9@        ������������������������       �                     @                                `f�<@r�q��?             2@                                `fF:@      �?             @        ������������������������       �                      @        ������������������������       �      �?             @        ������������������������       �                     (@                                   �?�����H�?            �F@                                   �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @               !                    4@��(\���?             D@                                    &@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        "       )                    �?г�wY;�?             A@       #       $                   �;@(;L]n�?             >@        ������������������������       �        	             .@        %       &                   �'@��S�ۿ?
             .@       ������������������������       �                     (@        '       (                    =@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        +       ^                 `f^@�������?4            �V@       ,       ?                   �E@�~�4_��?3             V@        -       >                    �?h+�v:�?             A@       .       /                 `fF)@����e��?            �@@        ������������������������       �                     @        0       1                   �@@|��?���?             ;@        ������������������������       �                      @        2       3                    �?� �	��?             9@        ������������������������       �                     �?        4       ;                    �?r�q��?             8@       5       6                     �?��.k���?             1@        ������������������������       �                     @        7       8                   @A@և���X�?             ,@        ������������������������       ��q�q�?             @        9       :                   @C@      �?              @        ������������������������       �                     @        ������������������������       ����Q��?             @        <       =                 03U@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        @       O                   �H@�����H�?             K@        A       D                    �?�㙢�c�?             7@        B       C                   �G@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        E       N                   �G@�����H�?             2@       F       M                    �?�IєX�?
             1@       G       L                     �?�8��8��?             (@       H       K                    G@      �?              @       I       J                 `f?@      �?             @       ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        P       U                    �?`Jj��?             ?@        Q       T                 ���Q@r�q��?             @       R       S                   �L@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        V       ]                    �?`2U0*��?             9@       W       X                   �N@���7�?             6@       ������������������������       �        
             2@        Y       \                 `f�2@      �?             @       Z       [                   �P@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        `       g                    �?������?1            �R@       a       b                    �?�Ń��̧?             E@       ������������������������       �                     6@        c       d                 ���`@P���Q�?             4@       ������������������������       �        	             0@        e       f                 Ъ�c@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        h       �                    @4���C�?            �@@       i       |                     �?`՟�G��?             ?@       j       s                    �?���Q��?             .@        k       l                    3@      �?              @        ������������������������       �                     �?        m       r                    �?؇���X�?             @       n       o                    >@r�q��?             @        ������������������������       �                     @        p       q                 �;�p@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        t       {                     @և���X�?             @       u       v                    F@�q�q�?             @        ������������������������       �                     @        w       x                 `f�R@�q�q�?             @        ������������������������       �                     �?        y       z                 03�S@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        }       �                    �?      �?	             0@       ~                          �3@��S���?             .@        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �                        ��Y7@x%[VY[�?�            �x@       �       �                    �?���f+�?�            `u@        �       �                    @f���M�?;            @W@       �       �                 ��.@��|�	��?9            �V@       �       �                    �?T�iA�?-            �Q@       �       �                 P��+@<��¤�?+             Q@       �       �                    1@�BE����?'             O@        �       �                    @�����H�?             "@        �       �                 P��%@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                 @3�@䯦s#�?!            �J@       �       �                    �?¦	^_�?             ?@        �       �                    7@8�Z$���?
             *@        ������������������������       �                     �?        �       �                 ���@�8��8��?	             (@        �       �                 0��@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@        �       �                   �;@b�2�tk�?
             2@       �       �                 �&B@d}h���?             ,@       �       �                 ���@      �?              @        ������������������������       �                      @        �       �                    4@      �?             @        ������������������������       �                      @        �       �                   �7@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 `�X!@      �?             6@        ������������������������       �                     @        �       �                 ��i#@     ��?
             0@        �       �                    �?�����H�?             "@       �       �                   �;@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?և���X�?             @       �       �                  �#@z�G�z�?             @       ������������������������       �                     @        �       �                    4@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                    ;@�����?             5@        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     .@        ������������������������       �                      @        �       �                    ,@� ��?�             o@        �       �                   X1@����X�?             @        ������������������������       �                     @        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �                         @@@��2(&�?�            @n@       �                        �v6@ZՏ�m|�?�            �h@       �                       ��i @��5�W�?             h@       �       �                   �0@u�����?_            �b@        ������������������������       �      �?             @        �       �                    �?д>��C�?]             b@       �       �                    �?� y���?U            �`@        �       �                    5@ףp=
�?             4@        �       �                 �{@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �:@�X�<ݺ?
             2@        ������������������������       �                      @        �       �                 ���@      �?             0@        ������������������������       �                     @        �       �                    =@�C��2(�?             &@       �       �                   @@ףp=
�?             $@       ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �<@�k�'7��?I            �\@       �       �                   �;@�+�ԗ�?@            �X@       �       �                    �?���B���?"             J@        ������������������������       �                      @        �       �                 ��L@z�G�z�?!             I@        �       �                   �:@�q�q�?             ;@       �       �                 �?$@��<b���?             7@       �       �                 ���@�t����?             1@        �       �                 �&b@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@        �       �                   �6@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                 @3�@�nkK�?             7@        ������������������������       �                     "@        �       �                   �3@@4և���?	             ,@        ������������������������       �      �?              @        ������������������������       �                     (@        �       �                    �?�q��/��?             G@        ������������������������       �        
             ,@        �       �                 ��) @     ��?             @@       �       �                  sW@ 	��p�?             =@        �       �                 pf�@      �?              @        ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                     5@        ������������������������       �                     @        �       �                    �?     ��?	             0@        ������������������������       �                     @        �       �                   �?@8�Z$���?             *@        ������������������������       �                     @        �       �                   �@�q�q�?             @        ������������������������       �                     �?        �       �                 �?�@z�G�z�?             @        ������������������������       �                     @        ������������������������       �      �?              @        �                          �?���!pc�?             &@       �       �                    3@�z�G��?             $@        ������������������������       �                     @        �                         �:@և���X�?             @       �                           5@      �?             @        ������������������������       �                      @                              ��@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?                                 �?���7�?              F@                                9@@4և���?             <@       ������������������������       �                     0@        	                      �̤0@r�q��?             (@       
                      ���"@�C��2(�?             &@        ������������������������       �                     @                                 (@z�G�z�?             @                               �<@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     0@        ������������������������       �                     @                                 �?��<b�ƥ?             G@        ������������������������       �                     @                                 �?��Y��]�?            �D@                                �?�?�|�?            �B@                               @F@�g�y��?             ?@                               �E@��S�ۿ?             .@       ������������������������       �                     (@                              @3�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     0@        ������������������������       �                     @        ������������������������       �                     @        !      &                   �?l�b�G��?!            �L@        "      #                �T)D@      �?             @        ������������������������       �                      @        $      %                   ;@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        '      (                   @���J��?            �I@        ������������������������       �                     3@        )      0                   @      �?             @@       *      +                   �?P���Q�?	             4@        ������������������������       �                     @        ,      -                ��T?@$�q-�?             *@       ������������������������       �                      @        .      /                   �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        �t�bh�h*h-K ��h/��R�(KM1KK��h]�B       P|@     0p@     �c@     �c@      a@     �Y@      �?     �Q@              O@      �?      "@      �?      @      �?                      @              @     �`@      ?@     �P@      $@      :@      @      @       @      @       @      @                       @      �?              6@      @      @              .@      @      @      @       @              �?      @      (@              D@      @      @       @               @      @             �B@      @      @       @               @      @             �@@      �?      =@      �?      .@              ,@      �?      (@               @      �?              �?       @              @             @Q@      5@     @Q@      3@      5@      *@      4@      *@      @              ,@      *@               @      ,@      &@      �?              *@      &@       @      "@              @       @      @       @      @      @       @      @              @       @      @       @      @                       @      �?              H@      @      3@      @      @       @      @                       @      0@       @      0@      �?      &@      �?      @      �?      @      �?      �?      �?       @              @              @              @                      �?      =@       @      @      �?       @      �?              �?       @              @              8@      �?      5@      �?      2@              @      �?       @      �?              �?       @              �?              @                       @      4@     �K@      �?     �D@              6@      �?      3@              0@      �?      @      �?                      @      3@      ,@      1@      ,@      "@      @      @       @              �?      @      �?      @      �?      @              �?      �?      �?                      �?      �?              @      @       @      @              @       @      �?      �?              �?      �?              �?      �?              �?               @       @       @      @              @       @                      �?       @             �r@     �Y@     �n@     �X@     �@@      N@      ?@      N@      =@     �D@      ;@     �D@      5@     �D@      �?       @      �?      �?      �?                      �?              @      4@     �@@      "@      6@       @      &@      �?              �?      &@      �?       @               @      �?                      "@      @      &@      @      &@      @      @               @      @      @       @              �?      @              @      �?                      @      @              &@      &@      @              @      &@      �?       @      �?      @      �?                      @               @      @      @      @      �?      @              �?      �?              �?      �?                       @      @               @               @      3@       @      @       @                      @              .@       @             `j@      C@       @      @              @       @      �?       @                      �?      j@     �@@     �d@      @@     �d@      =@     �^@      ;@       @       @      ^@      9@      \@      6@      2@       @      �?      �?      �?                      �?      1@      �?       @              .@      �?      @              $@      �?      "@      �?      @      �?       @              �?             �W@      4@     �T@      .@      E@      $@       @              D@      $@      2@      "@      2@      @      .@       @      @       @      @                       @      "@              @      @              @      @                      @      6@      �?      "@              *@      �?      �?      �?      (@             �D@      @      ,@              ;@      @      ;@       @      @       @      @              �?       @      5@                      @      &@      @              @      &@       @      @              @       @              �?      @      �?      @              �?      �?       @      @      @      @      @              @      @      �?      @               @      �?      �?      �?                      �?      @              �?              E@       @      :@       @      0@              $@       @      $@      �?      @              @      �?      @      �?      @                      �?      �?                      �?      0@                      @     �F@      �?      @              D@      �?      B@      �?      >@      �?      ,@      �?      (@               @      �?              �?       @              0@              @              @             �J@      @      @      @       @              �?      @              @      �?              I@      �?      3@              ?@      �?      3@      �?      @              (@      �?       @              @      �?              �?      @              (@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ:d�hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B�G         b                     @���x�W�?�           @�@                                   �?��$p�w�?�            �r@                                   �?��.N"Ҭ?U            @a@                                ��A@��p\�?            �D@                                `v7<@���!pc�?             &@       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     >@        	       
                    �?�a�O�?<            @X@       ������������������������       �        "             K@                                   6@ qP��B�?            �E@                                   �?      �?             @                                 �<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                    �C@               E                     �?�����?e            �c@              "                    �?�!>�R�?3            �T@               !                 �̾w@X�<ݚ�?             ;@                                 �1@�q�����?             9@        ������������������������       �                     @                                   �?և���X�?             5@                                  �?���|���?             &@        ������������������������       �                     @        ������������������������       �                     @                                ��+T@      �?             $@        ������������������������       �                      @                                ��hU@      �?              @        ������������������������       �                     @                                 @�pX@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        #       0                   �>@Dc}h��?#             L@        $       '                   �A@      �?             4@        %       &                   �;@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        (       -                    K@�	j*D�?             *@       )       ,                    H@�����H�?             "@       *       +                 03k:@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     @        .       /                 `fF<@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        1       D                    @tk~X��?             B@       2       =                  D0T@     ��?             @@       3       4                    �?���}<S�?             7@        ������������������������       �                     $@        5       <                   @K@8�Z$���?             *@        6       ;                    �?����X�?             @       7       8                 `fFJ@r�q��?             @        ������������������������       �                      @        9       :                    7@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        >       ?                   �D@X�<ݚ�?             "@        ������������������������       �                     @        @       A                   �G@z�G�z�?             @        ������������������������       �                     @        B       C                     @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        F       W                    �?�=A�F�?2             S@       G       H                    !@ i���t�?             �H@        ������������������������       �                     �?        I       V                 `��,@�8��8��?             H@       J       U                 ��\+@������?            �D@       K       R                    @@��(\���?             D@       L       Q                    5@ ��WV�?             :@        M       N                   �2@�C��2(�?             &@       ������������������������       �                     @        O       P                   �'@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �        
             .@        S       T                   �A@؇���X�?             ,@        ������������������������       ����Q��?             @        ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     @        X       _                    �?��}*_��?             ;@       Y       ^                   �@@��S�ۿ?
             .@        Z       [                    �?؇���X�?             @        ������������������������       �                     @        \       ]                   �H@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        `       a                    6@      �?             (@       ������������������������       �                     "@        ������������������������       �                     @        c       p                    @�g���l�?           �y@        d       e                    @�q�q�?             >@        ������������������������       �                     .@        f       g                    �?�q�q�?
             .@        ������������������������       �                     @        h       m                    �?X�<ݚ�?             "@       i       j                    @      �?             @        ������������������������       �                      @        k       l                    @      �?             @        ������������������������       �                     @        ������������������������       �                     �?        n       o                 ��T?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        q                          �?r^fx���?�            x@       r       �                    �?nb<��?�            Pu@        s       �                    �?�^�X�?>            @X@        t       �                    �?�4F����?            �D@        u       �                    �?��S���?
             .@       v       {                    5@���|���?             &@        w       z                    �?�q�q�?             @       x       y                    .@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        |       }                    :@      �?              @        ������������������������       �                     �?        ~       �                   �<@����X�?             @              �                    �?�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �7@�θ�?             :@        �       �                    �?      �?              @        �       �                   �0@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                 ��&@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                 ���@�����H�?             2@        ������������������������       �                      @        �       �                 �� @z�G�z�?	             $@       �       �                   @@�<ݚ�?             "@        ������������������������       �      �?             @        �       �                   �<@z�G�z�?             @        ������������������������       �                      @        �       �                    ?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                    1@Dc}h��?"             L@        ������������������������       �                     @        �       �                   �=@      �?              J@       �       �                    �?�7����?            �G@       �       �                    �?����>�?            �B@       �       �                 ���@�\��N��?             3@        ������������������������       �                     @        �       �                 ���@     ��?             0@        ������������������������       �                     @        �       �                    9@��
ц��?	             *@        ������������������������       �                     �?        �       �                    �?�q�q�?             (@       �       �                 pF @      �?             $@       �       �                 �&B@X�<ݚ�?             "@       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �8@�X�<ݺ?             2@        ������������������������       �                     �?        �       �                 03�@�IєX�?             1@        ������������������������       �                     @        �       �                 ��(@�C��2(�?             &@       ������������������������       �r�q��?             @        ������������������������       �                     @        �       �                 03�3@�z�G��?             $@       �       �                    �?և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �                          @yٯ���?�            �n@       �       �                    �?�֪u�_�?�            �m@       �       �                    �?T���ʴ�?            �h@       �       �                    O@�r&��K�?y            `g@       �       �                    �?\[j��?x             g@        �       �                   �@�q�����?             9@        �       �                   �3@      �?              @        �       �                 P��@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    4@�t����?             1@        ������������������������       �                     �?        �       �                   �9@      �?             0@        ������������������������       �                     @        �       �                   &@X�<ݚ�?             "@       �       �                 @3�@      �?              @        �       �                 �?�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ��� @z�G�z�?             @        ������������������������       �                     @        �       �                  SE"@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 �T�C@p=
ףp�?f             d@       �       �                   �0@ ��Ou��?b            �c@        �       �                 pf�@����X�?             @        ������������������������       �                     �?        �       �                 �̌!@�q�q�?             @       ������������������������       ����Q��?             @        ������������������������       �                     �?        �       �                 ���"@p���?^            �b@       �       �                   �>@�M8��p�?V             a@       �       �                   �8@��<b�ƥ?8             W@        ������������������������       �                    �C@        �       �                   �9@�&=�w��?            �J@        �       �                 @33@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �?$@`Ql�R�?            �G@        �       �                    =@؇���X�?             @       �       �                 pf�@z�G�z�?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     D@        �       �                   @@@�:�^���?            �F@        �       �                 �?�@X�<ݚ�?             "@        ������������������������       �                     @        �       �                 ��i @z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     B@        �       �                 ���#@r�q��?             (@        �       �                   �<@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                 pff0@�q�q�?             (@       �       �                    �?�z�G��?             $@       �       �                   @A@�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �                         @A@���@��?            �B@       �                         �9@�חF�P�?             ?@        �                       03#,@�z�G��?             $@       �       �                    3@      �?             @        ������������������������       �                      @                               ��@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                                 �?�����?             5@                                �?�����H�?             2@                                �>@      �?              @                               �.@؇���X�?             @        ������������������������       �                     @        	      
                   ;@      �?             @        ������������������������       �                      @                                 4@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     @                                 �?      �?             @                               �*@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @                                 @t��ճC�?             F@                                 �?H%u��?             9@                                 �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @                                �>@P���Q�?
             4@       ������������������������       �        	             3@        ������������������������       �                     �?        ������������������������       �                     3@        �t�bh�h*h-K ��h/��R�(KMKK��h]�B�       P{@     0q@      ]@     �f@      @     �`@      @      C@      @       @               @      @                      >@      �?      X@              K@      �?      E@      �?      @      �?      �?      �?                      �?               @             �C@      \@     �G@     �I@      @@      (@      .@      (@      *@              @      (@      "@      @      @              @      @              @      @               @      @      @      @               @      @              @       @                       @     �C@      1@      $@      $@      @      �?              �?      @              @      "@      �?       @      �?      @              �?      �?       @              @      @      �?      @                      �?      =@      @      9@      @      5@       @      $@              &@       @      @       @      @      �?       @              @      �?      @                      �?              �?      @              @      @              @      @      �?      @              �?      �?              �?      �?              @             �N@      .@      F@      @              �?      F@      @     �B@      @     �B@      @      9@      �?      $@      �?      @              @      �?       @      �?      �?              .@              (@       @      @       @      "@                      �?      @              1@      $@      ,@      �?      @      �?      @               @      �?              �?       @               @              @      "@              "@      @             t@     �W@      $@      4@              .@      $@      @      @              @      @      @      @       @              �?      @              @      �?              �?       @      �?                       @     ps@     �R@     �p@     �Q@     �P@      >@      <@      *@       @      @      @      @       @      �?      �?      �?              �?      �?              �?               @      @              �?       @      @       @      @              @       @                      �?      @              4@      @      @      @       @       @       @                       @       @       @       @                       @      0@       @       @               @       @      @       @      @      �?      @      �?       @               @      �?              �?       @              �?             �C@      1@              @     �C@      *@      A@      *@      ;@      $@      $@      "@      @              @      "@              @      @      @              �?      @      @      @      @      @      @      @      @              �?      �?               @              1@      �?      �?              0@      �?      @              $@      �?      @      �?      @              @      @      @      @              @      @              @              @             `i@     �D@     `h@     �D@     �d@     �@@     �c@      <@     �c@      :@      *@      (@      �?      @      �?       @               @      �?                      @      (@      @              �?      (@      @      @              @      @      @      @      �?       @      �?                       @      @      �?      @              �?      �?              �?      �?                      �?     @b@      ,@     @b@      $@      @       @      �?              @       @      @       @      �?             �a@       @     ``@      @     �V@       @     �C@             �I@       @      @      �?              �?      @              G@      �?      @      �?      @      �?       @               @      �?       @              D@             �D@      @      @      @      @              �?      @              @      �?              B@              $@       @      @       @      @                       @      @                      @               @      @      @      @      @      @      @              @      @              �?                       @      =@       @      :@      @      @      @      @      @       @              �?      @      �?                      @      @              3@       @      0@       @      @       @      @      �?      @              @      �?       @              �?      �?              �?      �?                      �?      $@              @              @      @      �?      @      �?                      @       @               @             �D@      @      6@      @      @       @      @                       @      3@      �?      3@                      �?      3@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�I]fhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtK�huh*h-K ��h/��R�(KK�h|�B�<         N                 `f�%@������?�           @�@                                   �?��U'�?�            �q@                                pF @Np�����?"            �I@                                  �?����X�?             <@              
                 ���@@�0�!��?             1@               	                 �Y�@      �?             @                               03�@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        	             *@                                   0@�eP*L��?	             &@        ������������������������       �                      @                                   8@�q�q�?             "@        ������������������������       �                     @                                   �?���Q��?             @                               �?�@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?                                    @��<b���?             7@        ������������������������       �                     @                                   3@�}�+r��?
             3@        ������������������������       �                     �?        ������������������������       �        	             2@                                ���@$]^z���?�             m@        ������������������������       �                     9@               1                    �?�����H�?�            �i@               0                    �?<ݚ)�?             B@                                  9@r٣����?            �@@        ������������������������       �                     @                /                   �=@r�q��?             >@       !       "                 ���@�E��ӭ�?             2@        ������������������������       �                     @        #       .                    �?X�Cc�?             ,@       $       +                 03s@�n_Y�K�?             *@       %       *                   @<@���|���?	             &@       &       '                    �?���Q��?             $@        ������������������������       �      �?              @        (       )                 ��(@      �?              @       ������������������������       �և���X�?             @        ������������������������       �                     �?        ������������������������       �                     �?        ,       -                   �<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                     @        2       G                   @C@l�b�G��?h            `e@       3       4                 ��@F��}��?Y            @b@        ������������������������       �                     @        5       D                    $@��K˱F�?X            �a@       6       C                    �?�z�N��?Q            ``@       7       8                 �?�@�U���?P            �_@        ������������������������       �        &            �P@        9       >                 @3�@�.ߴ#�?*            �N@        :       ;                    >@"pc�
�?             &@        ������������������������       �                     @        <       =                    �?����X�?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ?       B                 ��Y @p���?$             I@       @       A                   �3@h�����?             <@        ������������������������       �      �?              @        ������������������������       �                     :@        ������������������������       �                     6@        ������������������������       �                     @        E       F                   �5@r�q��?             (@        ������������������������       ����Q��?             @        ������������������������       �                     @        H       I                 �?�@�J�4�?             9@       ������������������������       �                     *@        J       M                    �?�q�q�?             (@       K       L                 @3�@���Q��?             $@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        O       �                    @��ߚ���?           �z@       P       {                    �?��^@=��?�            �x@        Q       ^                     @B�#-g�?r            �g@       R       S                    @��.N"Ҭ?U            @a@        ������������������������       �                     @        T       ]                     �?���б�?T            �`@       U       V                    �?`׀�:M�?/            �R@       ������������������������       �        (             O@        W       X                   �8@�8��8��?             (@       ������������������������       �                      @        Y       Z                    �?      �?             @        ������������������������       �                      @        [       \                 ���`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        %            �N@        _       d                   �6@�F�j��?            �J@        `       c                   �"@      �?             0@        a       b                 �>1@X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        e       z                 `v�6@�Gi����?            �B@       f       y                    @     ��?             @@       g       h                   �;@�4�����?             ?@        ������������������������       �                     @        i       v                    �?��}*_��?             ;@       j       u                   �D@�X����?             6@       k       p                 pF�-@����X�?
             5@        l       m                    �?z�G�z�?             @        ������������������������       �                      @        n       o                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        q       r                   �=@      �?             0@       ������������������������       �                     $@        s       t                   �@@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        w       x                   �<@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        |       �                    �?�h0����?            @i@       }       �                 �ܵ<@�=A�F�?_             c@       ~                          �9@�Ra����?9             V@        ������������������������       �                     4@        �       �                   �:@��hJ,�?-             Q@        �       �                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�? Da�?+            �O@       �       �                     @X��Oԣ�?*             O@       �       �                    �?�T|n�q�?            �E@        ������������������������       �                     @        �       �                     �?:�&���?            �C@        �       �                 03k:@8�Z$���?	             *@        �       �                   �A@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    J@�C��2(�?             &@        �       �                   @G@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 `f�)@���B���?             :@        ������������������������       �                      @        �       �                   �;@�q�q�?             8@        ������������������������       �                     @        �       �                   �@@�d�����?             3@        �       �                    �?      �?             @        ������������������������       �                     �?        �       �                   �7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    F@�r����?             .@       �       �                    �?z�G�z�?             $@       �       �                    C@���Q��?             @       ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     3@        ������������������������       �                     �?        �       �                     @     ��?&             P@       �       �                     �?������?#             N@       �       �                   �>@�c�Α�?!             M@        �       �                 ���=@�q�q�?             "@        �       �                   �E@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �J@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                 ��9L@�����?            �H@       �       �                    �?�8��8��?             8@       �       �                   �I@      �?
             0@       �       �                    �?@4և���?             ,@        ������������������������       �                     @        �       �                   �=@�C��2(�?             &@       �       �                 ��yC@؇���X�?             @        �       �                   �@@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   @A@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   @G@`�Q��?             9@       �       �                   �;@��+7��?
             7@        �       �                    �?�q�q�?             @        ������������������������       �                     @        �       �                   �5@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?�t����?             1@        ������������������������       �                     �?        �       �                   �@@      �?             0@        �       �                    �?r�q��?             @        ������������������������       �                      @        �       �                    >@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?z�):���?              I@        �       �                      @      �?              @       �       �                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �3@�G��l��?             E@        �       �                    �?     ��?             0@        �       �                 ���*@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        �       �                    �?$��m��?             :@        �       �                    )@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    (@���Q��?             4@        ������������������������       �                     @        �       �                     �?؇���X�?
             ,@        �       �                     @      �?              @       �       �                    F@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @������?             B@        �       �                    �?�8��8��?             (@        ������������������������       �                     @        �       �                    @z�G�z�?             @       �       �                    @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     8@        �t�b��      h�h*h-K ��h/��R�(KK�KK��h]�B0        |@     `p@     `m@      H@      :@      9@       @      4@      @      ,@      @      �?      �?      �?      �?                      �?       @                      *@      @      @       @              @      @              @      @       @       @       @       @                       @      �?              2@      @              @      2@      �?              �?      2@              j@      7@      9@              g@      7@      9@      &@      9@       @              @      9@      @      *@      @      @              "@      @       @      @      @      @      @      @      �?      �?      @      @      @      @      �?              �?              �?      �?      �?                      �?      �?              (@                      @     �c@      (@     @a@       @              @     @a@      @      `@      @      _@      @     �P@              M@      @      "@       @      @              @       @      @       @      �?             �H@      �?      ;@      �?      �?      �?      :@              6@              @              $@       @      @       @      @              5@      @      *@               @      @      @      @              @      @               @             �j@     �j@     �f@     �j@      ?@      d@      @     �`@      @              �?     �`@      �?     @R@              O@      �?      &@               @      �?      @               @      �?      �?              �?      �?                     �N@      ;@      :@      (@      @      @      @              @      @              @              .@      6@      $@      6@      $@      5@              @      $@      1@      @      .@      @      .@      @      �?       @               @      �?              �?       @               @      ,@              $@       @      @       @                      @      �?              @       @      @                       @              �?      @             �b@     �J@     �^@      >@     �S@      $@      4@              M@      $@      @       @               @      @             �K@       @     �K@      @      B@      @      @              @@      @      &@       @      �?      �?      �?                      �?      $@      �?      @      �?      @                      �?      @              5@      @       @              3@      @      @              ,@      @      �?      @              �?      �?       @      �?                       @      *@       @       @       @      @       @      @      �?              �?      @              @              3@                      �?      F@      4@      F@      0@      E@      0@      @      @      �?      �?              �?      �?               @      @              @       @             �C@      $@      6@       @      ,@       @      *@      �?      @              $@      �?      @      �?      �?      �?      �?                      �?      @              @              �?      �?      �?                      �?       @              1@       @      1@      @       @      @              @       @      �?       @                      �?      .@       @              �?      .@      �?      @      �?       @              @      �?      @                      �?      $@                       @       @                      @      ;@      7@      @      �?      @      �?      @                      �?      @              4@      6@      @      *@      @      �?              �?      @                      (@      1@      "@      @      �?              �?      @              (@       @              @      (@       @      @       @      @       @               @      @              �?              @             �A@      �?      &@      �?      @              @      �?       @      �?       @                      �?       @              8@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�޵#hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMKhuh*h-K ��h/��R�(KMK��h|�B�R                         `f~I@~�Я��?�           @�@              �                    �?��}y.��?e           ȁ@              �                    @�5�l	�?           0|@              ;                    �?��n����?           �{@                                ��Y@z)�J'c�?G            @]@        ������������������������       �                     @                                    @�{���2�?C            �[@                                `��,@�5��?             ;@        	       
                    �?؇���X�?             @       ������������������������       �                     @                                  @E@      �?             @        ������������������������       �                     @        ������������������������       �                     �?                                   E@      �?             4@                                  �?�r����?             .@       ������������������������       �                     *@        ������������������������       �                      @                                  �L@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @                                  �0@\`*�s�?3             U@                                �y.@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?               $                    �?��مD�?.            @S@                                  �7@�J�4�?             9@                                  �3@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   ;@�LQ�1	�?             7@        ������������������������       �                     @                #                    �?R���Q�?             4@       !       "                    �?�S����?             3@        ������������������������       �                     @        ������������������������       �        	             0@        ������������������������       �                     �?        %       4                 03�'@      �?             J@       &       3                    >@>A�F<�?             C@       '       (                 ��@H�V�e��?             A@        ������������������������       �                     @        )       0                    �?������?             ;@        *       /                 `f�@��
ц��?             *@       +       ,                   �8@�q�q�?             "@        ������������������������       �                     �?        -       .                 ���@      �?              @        ������������������������       �                     �?        ������������������������       �����X�?             @        ������������������������       �                     @        1       2                   �<@@4և���?	             ,@       ������������������������       �                     *@        ������������������������       �                     �?        ������������������������       �                     @        5       :                 03�7@և���X�?             ,@       6       9                   `3@      �?              @       7       8                    �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        <       �                   �R@�GN�z�?�            �t@       =       t                     @DV��%�?�            �t@        >       C                    �?*AA,�P�?G            @^@        ?       B                  �v7@z�G�z�?             9@       @       A                   �;@�E��ӭ�?
             2@        ������������������������       �                     @        ������������������������       �                     *@        ������������������������       �                     @        D       K                   �;@     ��?7             X@        E       J                    5@���N8�?             5@        F       G                   �1@�����H�?             "@        ������������������������       �                      @        H       I                   �'@؇���X�?             @       ������������������������       �r�q��?             @        ������������������������       �                     �?        ������������������������       �                     (@        L       s                    �?��n�?,            �R@       M       f                   �B@H�V�e��?(             Q@       N       O                 `fF)@��Hg���?            �F@        ������������������������       �                     (@        P       e                 `f�D@�q�q�?            �@@       Q       `                    @@��>4և�?             <@       R       _                   �A@�����?             3@       S       ^                   �<@�E��ӭ�?
             2@       T       [                     �?     ��?             0@       U       V                 `fF:@�	j*D�?             *@        ������������������������       �                     @        W       Z                   �>@���Q��?             $@       X       Y                 `f�<@      �?              @       ������������������������       �և���X�?             @        ������������������������       �                     �?        ������������������������       �                      @        \       ]                   �*@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        a       d                 ��$:@X�<ݚ�?             "@       b       c                   @A@և���X�?             @       ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        g       h                   `G@�LQ�1	�?             7@        ������������������������       �                     "@        i       n                     �?d}h���?	             ,@        j       m                 `f�<@r�q��?             @       k       l                    K@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        o       p                   @N@      �?              @       ������������������������       �                     @        q       r                   �P@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        u       �                 @3�@ԩ��/�?�            �i@       v       �                   @@@������?J            �]@       w       �                 �?�@Nṧ'
�?:            �W@       x       �                    �?�A+K&:�?1             S@        y       z                    4@X�<ݚ�?             "@        ������������������������       �                      @        {       �                   �@����X�?             @       |       �                 �&B@r�q��?             @       }       ~                 ��@      �?             @        ������������������������       �                     �?               �                   �7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                 ��@�Y����?*            �P@        �       �                 ��@և���X�?             @       �       �                    6@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                 �{@�r����?&             N@       �       �                 �?$@z�G�z�?             D@       �       �                    7@@4և���?             <@        ������������������������       �        	             1@        �       �                 ���@"pc�
�?
             &@        �       �                 �&b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    ;@�����H�?             "@        ������������������������       �                      @        �       �                    =@؇���X�?             @       �       �                 pf�@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ��L@      �?             (@        �       �                   �8@���Q��?             @       �       �                   �5@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    :@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     4@        �       �                   �9@�\��N��?	             3@        �       �                   �4@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?z�G�z�?             $@        ������������������������       �                     @        �       �                   �?@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �C@ �q�q�?             8@        �       �                 �?�@ףp=
�?             $@       ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        	             ,@        �       �                 ���"@�Ra����?>             V@       �       �                    �?�X�<ݺ?$             K@        ������������������������       �                     @        �       �                   �0@=QcG��?             �G@        ������������������������       �      �?             @        �       �                 ��i @ qP��B�?            �E@       �       �                    ?@h�����?             <@       ������������������������       �                     1@        �       �                   �@@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �        
             .@        �       �                 0S�*@H�V�e��?             A@        �       �                    3@�q�q�?	             (@        ������������������������       �                      @        �       �                    �?�z�G��?             $@       �       �                   �<@      �?              @        ������������������������       �                     @        �       �                   �@@      �?             @        ������������������������       �                      @        �       �                    I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�C��2(�?             6@        �       �                   �=@�q�q�?             @       �       �                    5@      �?             @        ������������������������       �                     �?        �       �                    9@�q�q�?             @        ������������������������       �                     �?        �       �                    ;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     0@        ������������������������       �                      @        ������������������������       �                     @        �       �                 ��97@�m����?L            �]@        �       �                 P�@�2�o�U�?!            �K@        ������������������������       �                      @        �       �                 @�+@�#ʆA��?             �J@        ������������������������       �                     ,@        �       �                    @�n_Y�K�?            �C@       �       �                     @^H���+�?            �B@        ������������������������       �                      @        �       �                 ���.@П[;U��?             =@        �       �                   �<@�<ݚ�?             "@        ������������������������       �                     @        �       �                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    3@�z�G��?             4@       �       �                    �?      �?             $@       �       �                     @����X�?             @        �       �                    +@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 pff0@ףp=
�?             $@        �       �                 �y�/@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?���h%��?+            �O@       �       �                 м�9@     ��?             @@        ������������������������       �                     @        �       �                 03;@��
ц��?             :@        ������������������������       �                      @        �       �                     @�q�q�?             2@        ������������������������       �                     @        �       �                    @؇���X�?
             ,@        �       �                 ��T?@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@                                  @�n`���?             ?@                                �C@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @                                  @HP�s��?             9@                                 �?8�Z$���?             *@        ������������������������       �                     @                                  @�<ݚ�?             "@             	                   �?�q�q�?             @        ������������������������       �                     �?        
                        �B@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        	             (@                                 �?OX���?W            �a@                                �?���Lͩ�?-            �R@        ������������������������       �                     7@                                �<@���c���?             J@                                �8@R�}e�.�?             :@                                 @@4և���?             ,@        ������������������������       �                     �?        ������������������������       �                     *@                                 �?      �?             (@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     :@              F                  @I@�ʻ����?*             Q@             A                   �?��k��?$            �J@             .                   �?X��ʑ��?            �E@                                �8@X�<ݚ�?             2@        ������������������������       �                     @               '                   �?�q�q�?
             .@        !      &                   �?���Q��?             @       "      #                  �?@      �?             @        ������������������������       �                      @        $      %                  @D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        (      -                p"�X@z�G�z�?             $@       )      ,                   C@�����H�?             "@       *      +                  �:@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        /      >                    @�q�����?             9@       0      =                    �?���Q��?             4@       1      <                ���[@��.k���?             1@       2      ;                  �C@X�Cc�?             ,@       3      8                   �?      �?             $@       4      7                `f�N@      �?              @       5      6                `fFJ@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        9      :                   =@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ?      @                   >@z�G�z�?             @        ������������������������       �      �?              @        ������������������������       �                     @        B      E                     @�z�G��?             $@       C      D                �̰f@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        G      J                   �?��S�ۿ?             .@        H      I                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     *@        �t�bh�h*h-K ��h/��R�(KMKKK��h]�B�       �{@     �p@     �x@     `e@      u@     @\@      u@     @[@     �T@      A@      @             @S@      A@      0@      &@      �?      @              @      �?      @              @      �?              .@      @      *@       @      *@                       @       @      @              @       @             �N@      7@      �?      @              @      �?              N@      1@      5@      @      �?      �?      �?                      �?      4@      @      @              1@      @      0@      @              @      0@              �?             �C@      *@      ?@      @      ;@      @      @              4@      @      @      @      @      @      �?               @      @              �?       @      @      @              *@      �?      *@                      �?      @               @      @       @      @       @      @              @       @                      @      @             �o@     �R@     �o@     @R@     �U@     �A@      @      4@      @      *@      @                      *@              @     @T@      .@      4@      �?       @      �?       @              @      �?      @      �?      �?              (@             �N@      ,@      K@      ,@      A@      &@      (@              6@      &@      1@      &@      *@      @      *@      @      &@      @      "@      @      @              @      @      @      @      @      @              �?       @               @      �?              �?       @               @                      �?      @      @      @      @      @      @      �?                       @      @              4@      @      "@              &@      @      @      �?      @      �?              �?      @              �?              @       @      @              @       @               @      @              @              e@      C@     �V@      <@      Q@      ;@     �M@      1@      @      @       @               @      @      �?      @      �?      @              �?      �?       @               @      �?                       @      �?             �K@      (@      @      @      @       @      @                       @               @      J@       @      @@       @      :@       @      1@              "@       @      �?      �?      �?                      �?       @      �?       @              @      �?      @      �?      @                      �?      �?              @      @       @      @       @      �?              �?       @                       @      @      @      @                      @      4@              "@      $@      @       @               @      @               @       @              @       @       @               @       @              7@      �?      "@      �?      @               @      �?              �?       @              ,@             �S@      $@     �I@      @      @              F@      @       @       @      E@      �?      ;@      �?      1@              $@      �?              �?      $@              .@              ;@      @      @      @               @      @      @      @      @      @              �?      @               @      �?      �?      �?                      �?       @              4@       @      @       @       @       @      �?              �?       @              �?      �?      �?      �?                      �?       @              0@                       @              @      N@      M@      1@      C@       @              .@      C@              ,@      .@      8@      *@      8@               @      *@      0@      @       @      @              @       @               @      @              @      ,@      @      @      @       @      �?       @               @      �?              @                      @      �?      "@      �?      �?              �?      �?                       @       @             �E@      4@      2@      ,@      @              (@      ,@               @      (@      @              @      (@       @      @       @      @                       @      "@              9@      @       @      @              @       @              7@       @      &@       @      @              @       @      @       @      �?              @       @               @      @              @              (@             �F@     �X@      @      Q@              7@      @     �F@      @      3@      �?      *@      �?                      *@      @      @              @      @                      :@      C@      >@      8@      =@      5@      6@       @      $@      @              @      $@      @       @      @      �?       @              �?      �?              �?      �?                      �?       @       @      �?       @      �?      @              @      �?                      @      �?              *@      (@      (@       @      "@       @      "@      @      @      @      @      @      �?      @      �?                      @      @              �?      �?      �?                      �?      @                      @      @              �?      @      �?      �?              @      @      @       @      @              @       @              �?              ,@      �?      �?      �?      �?                      �?      *@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�G�hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM;huh*h-K ��h/��R�(KM;��h|�B�N         ,                   �1@z����?�           @�@               	                     @d��0u��?:            �V@                                    �?      �?             @@        ������������������������       �                     $@                                   �?���7�?             6@                                  �&@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        
             3@        
                           @П[;U��?&             M@                                  #@�4�����?             ?@        ������������������������       �                     (@                                   �?�\��N��?             3@                                  �?���Q��?	             .@                                  �?�z�G��?             $@                                  (@      �?              @        ������������������������       �                     �?                                  �0@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?                                �&�)@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                �̌!@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @               +                    @�+$�jP�?             ;@                                  @      �?             4@        ������������������������       �                     @               $                    �?�t����?             1@                #                 ��T?@���Q��?             @       !       "                 ���3@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        %       *                    @r�q��?	             (@        &       '                    �?���Q��?             @        ������������������������       �                      @        (       )                    @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        -       �                     @f��yr}�?�           p�@        .       C                    �?.k����?�             q@        /       B                   �;@ ѯ��?F            �Z@        0       1                    �?�p ��?            �D@        ������������������������       �                     &@        2       =                    �?z�G�z�?             >@        3       4                     �?�q�q�?             (@        ������������������������       �                      @        5       :                   �9@���Q��?             $@       6       9                    �?r�q��?             @        7       8                   �6@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ;       <                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        >       ?                   �8@�����H�?	             2@       ������������������������       �                     .@        @       A                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        /            �P@        D       {                     �?��`���?c            �d@       E       J                    :@�5��
J�?5             W@        F       I                     @���Q��?             @       G       H                 8�T@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        K       Z                    �?&[i`��?2            �U@        L       Y                    �?r�q��?             8@       M       T                   @G@������?	             .@       N       S                    �?z�G�z�?             $@       O       R                   �?@����X�?             @       P       Q                 �ܵ<@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        U       X                 @�pX@���Q��?             @       V       W                 ��L@@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     "@        [       d                 `f�;@���N8�?%            �O@        \       ]                 ��$:@8�A�0��?             6@        ������������������������       �                     @        ^       _                 03k:@      �?	             2@        ������������������������       �                     @        `       c                   �J@X�Cc�?             ,@       a       b                   @B@����X�?             @        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     @        e       z                    R@�p ��?            �D@       f       y                    J@      �?             D@       g       v                    �?r�q��?             >@       h       u                    �?؇���X�?             <@       i       t                   �@@$�q-�?             :@       j       q                    >@r�q��?	             (@       k       l                   �@@�����H�?             "@        ������������������������       �                     @        m       p                    �?z�G�z�?             @       n       o                 ��yC@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        r       s                   @K@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     ,@        ������������������������       �                      @        w       x                 ���Y@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     �?        |       }                    �?F��}��?.            @R@        ������������������������       �                     ,@        ~       �                    �? ,��-�?'            �M@              �                   �<@��p\�?            �D@        �       �                   �'@�t����?             1@        ������������������������       �                     @        �       �                   �;@z�G�z�?             $@       ������������������������       �                     @        �       �                   �*@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   @D@ �q�q�?             8@       ������������������������       �                     .@        �       �                   �F@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�X�<ݺ?             2@       �       �                   �7@$�q-�?             *@        ������������������������       �                     @        �       �                   �:@�����H�?             "@       �       �                   �@@      �?              @        �       �                   �<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       2                  �@@���l��?�            �u@       �       1                   @������?�            �r@       �       .                   @��J��?�            @r@       �       !                  �?@@E>���?�            r@       �                       ��.@��v4Ք�?�            �p@       �       �                   �;@h�37*��?�            `k@       �       �                   �:@@��,*�?J            �]@       �       �                   �2@���@��?F            �[@        �       �                    �?�n_Y�K�?	             *@       �       �                    �?���Q��?             $@        �       �                 P��@z�G�z�?             @        ������������������������       �                      @        �       �                 ��!@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                 xF4!@�q�q�?             @        ������������������������       �                     �?        �       �                 ��'@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �@�[$�G�?=            �X@       �       �                    �?f�Sc��?            �H@        �       �                    8@z�G�z�?             .@       �       �                   �5@ףp=
�?             $@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                 �&B@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �3@@�0�!��?             A@        ������������������������       �                     @        �       �                    �?�n`���?             ?@       �       �                 �� @д>��C�?             =@        ������������������������       �                     �?        �       �                   �8@؇���X�?             <@       �       �                    7@"pc�
�?             6@       �       �                 03�@�S����?             3@        ������������������������       �                     @        �       �                 ���@z�G�z�?
             .@        ������������������������       �                     �?        �       �                    �?؇���X�?	             ,@        �       �                    5@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 @�@�C��2(�?             &@       ������������������������       �                     @        �       �                 ��L@z�G�z�?             @       �       �                   �5@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                   �@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                 �&B@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �3@@�E�x�?            �H@        �       �                 �?�@؇���X�?             @        ������������������������       �                     @        �       �                 `�8"@      �?             @        ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     E@        ������������������������       �                      @        �       �                    �?R���Q�?=             Y@        �       �                   �>@���|���?             6@       �       �                    =@�q�q�?             5@       �       �                  ��@��Q��?
             4@       �       �                    �?���|���?             &@       �       �                    �?�<ݚ�?             "@        ������������������������       �                     @        �       �                 �&B@�q�q�?             @       ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�:�^���?1            �S@        �       �                   @@     ��?	             0@       ������������������������       �                      @        �       �                 H�Z&@      �?              @       �       �                   �<@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �                          �?`Jj��?(             O@       �       �                    �?��S�ۿ?&             N@        �       �                 03�@���}<S�?             7@        ������������������������       �                     @        �       �                 ��(@      �?	             0@       �       �                   �<@؇���X�?             ,@       ������������������������       �                     $@        �       �                    >@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �                       ��) @@-�_ .�?            �B@       �                         �<@(;L]n�?             >@       �                       �?$@ �q�q�?             8@                               ��,@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     2@        ������������������������       �                     @                              pf� @؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        	                         �?����3��?#             J@        
                         ;@D�n�3�?             3@                              pff0@      �?              @        ������������������������       �                     �?        ������������������������       �                     @                              �T)D@�C��2(�?             &@       ������������������������       �                     @        ������������������������       �z�G�z�?             @                                 �?�q�q�?            �@@                                 �?�q�q�?             .@        ������������������������       �                     "@                                 �?r�q��?             @                                 ;@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                                �:@�X�<ݺ?             2@        ������������������������       �                     @                                  �?�C��2(�?             &@                                �?ףp=
�?             $@       ������������������������       �                      @                                 �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        "      -                  @@@      �?             2@       #      ,                �!B@�	j*D�?             *@       $      +                   �?���Q��?             $@       %      &                  �@      �?              @        ������������������������       �                      @        '      (                �?�@�q�q�?             @        ������������������������       �                     �?        )      *                @3�@z�G�z�?             @       ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        /      0                  �>@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        3      4                �?�@�NW���?             �J@       ������������������������       �                     <@        5      6                   �?�J�4�?             9@        ������������������������       �                     @        7      :                @3�@"pc�
�?             6@        8      9                  �D@z�G�z�?             @       ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �        
             1@        �t�bh�h*h-K ��h/��R�(KM;KK��h]�B�       �{@     �p@     �@@     �L@      �?      ?@              $@      �?      5@      �?       @      �?                       @              3@      @@      :@      $@      5@              (@      $@      "@      @      "@      @      @       @      @      �?              �?      @              @      �?              �?      �?              �?      �?              @       @               @      @              @              6@      @      .@      @      @              (@      @       @      @       @      �?              �?       @                       @      $@       @      @       @       @              �?       @      �?                       @      @              @             �y@      j@      b@     �_@      @     @Y@      @     �A@              &@      @      8@      @       @               @      @      @      �?      @      �?      �?              �?      �?                      @      @      �?              �?      @               @      0@              .@       @      �?              �?       @                     �P@     `a@      :@     �Q@      6@       @      @      �?      @              @      �?              �?              Q@      3@      4@      @      &@      @       @       @      @       @      @      �?      @                      �?              �?      @              @       @      �?       @      �?                       @       @              "@              H@      .@      *@      "@      @              "@      "@              @      "@      @       @      @       @       @              @      @             �A@      @     �A@      @      9@      @      8@      @      8@       @      $@       @       @      �?      @              @      �?      @      �?              �?      @              �?               @      �?       @                      �?      ,@                       @      �?      �?              �?      �?              $@                      �?     @Q@      @      ,@             �K@      @      C@      @      .@       @      @               @       @      @              @       @               @      @              7@      �?      .@               @      �?              �?       @              1@      �?      (@      �?      @               @      �?      @      �?      �?      �?      �?                      �?      @              �?              @             �p@     @T@     �k@     @S@     �j@     @S@     �j@     �R@     �i@     �P@     �e@     �G@     �U@      @@     �U@      8@       @      @      @      @      �?      @               @      �?       @      �?                       @      @               @      �?      �?              �?      �?              �?      �?             �S@      3@      ?@      2@      @      (@      �?      "@      �?      �?      �?                      �?               @       @      @       @                      @      <@      @      @              9@      @      8@      @              �?      8@      @      2@      @      0@      @      @              (@      @              �?      (@       @       @      �?              �?       @              $@      �?      @              @      �?       @      �?              �?       @               @               @      �?              �?       @              @              �?      �?              �?      �?              H@      �?      @      �?      @              @      �?      �?      �?       @              E@                       @     @U@      .@      ,@       @      ,@      @      *@      @      @      @       @      @              @       @      @       @      �?              @       @              "@              �?                      �?     �Q@      @      *@      @       @              @      @      @      @      @                      @       @              M@      @      L@      @      5@       @      @              ,@       @      (@       @      $@               @       @               @       @               @             �A@       @      =@      �?      7@      �?      @      �?      @                      �?      2@              @              @      �?              �?      @               @             �@@      3@      &@       @      �?      @      �?                      @      $@      �?      @              @      �?      6@      &@      @      $@              "@      @      �?       @      �?       @                      �?      @              1@      �?      @              $@      �?      "@      �?       @              �?      �?      �?                      �?      �?              "@      "@      @      "@      @      @       @      @               @       @      @      �?              �?      @      �?       @               @       @                      @      @              �?       @      �?                       @      @             �H@      @      <@              5@      @      @              2@      @      �?      @      �?       @               @      1@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ���JhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B@D         z                     @�VM�?�           @�@               W                    �?T �����?�             s@              <                     �?�3�w�?�             m@              3                 03?U@H������?J            @^@              
                    �?��C���?8            �W@               	                 03[=@�}�+r��?             3@                                `v7<@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        
             0@                                   �?������?+            �R@                                  �:@      �?
             4@        ������������������������       �                     @                                   ?@j���� �?	             1@                                  �?���!pc�?             &@                               ���<@�z�G��?             $@       ������������������������       �                     @                                03SA@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?                                ��>@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @                                  �;@"pc�
�?!            �K@                                `f�D@���Q��?             @        ������������������������       �                     �?                                   7@      �?             @        ������������������������       �                      @        ������������������������       �                      @               2                   @J@�:pΈ��?             I@               1                    �?��G���?            �B@       !       0                   �G@ �o_��?             9@       "       #                 ��I/@"pc�
�?             6@        ������������������������       �                      @        $       /                   �E@����X�?
             ,@       %       .                   �A@���|���?             &@       &       -                 ��yC@�z�G��?             $@       '       ,                   �A@      �?             @       (       +                   �<@      �?             @       )       *                   `@@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     (@        ������������������������       �                     *@        4       9                   �H@�<ݚ�?             ;@       5       6                 ���X@�LQ�1	�?             7@        ������������������������       �                     &@        7       8                    �?      �?
             (@       ������������������������       �                     "@        ������������������������       �                     @        :       ;                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        =       D                    �?����X�?@             \@        >       ?                   �2@h�����?             <@       ������������������������       �        
             3@        @       C                   �6@�����H�?             "@        A       B                   �<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        E       V                    �?(�s���?/             U@       F       S                   @N@$�q-�?&            @P@       G       H                   �;@�]0��<�?$            �N@        ������������������������       �                     7@        I       R                   �*@�}�+r��?             C@       J       K                 `fF)@�KM�]�?             3@        ������������������������       �                      @        L       M                    =@"pc�
�?	             &@        ������������������������       �                     �?        N       O                   @D@ףp=
�?             $@       ������������������������       �                     @        P       Q                   �F@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     3@        T       U                   �P@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             3@        X       i                     �?:PZ(8?�?,            @R@        Y       \                    �?�s��:��?             C@        Z       [                    '@��S�ۿ?
             .@        ������������������������       �                     �?        ������������������������       �        	             ,@        ]       h                 @�:x@8����?             7@       ^       g                 ��Ub@���!pc�?             6@       _       d                    �?      �?             0@       `       a                    �?      �?              @        ������������������������       �                     @        b       c                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        e       f                 03�S@      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        j       y                   �K@z�G�z�?            �A@       k       r                   @A@6YE�t�?            �@@       l       m                    �?���N8�?             5@        ������������������������       �                     @        n       o                    '@@4և���?
             ,@       ������������������������       �                      @        p       q                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        s       x                    �?�q�q�?             (@       t       u                    :@z�G�z�?             $@        ������������������������       �                     @        v       w                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        {       �                    �?���n�?�            `y@        |       �                    �?Hث3���?C            @]@        }       �                    �?r�q��?             E@       ~       �                    �?�'�`d�?            �@@               �                    :@�C��2(�?             &@        ������������������������       �                     @        �       �                 ��y&@      �?              @        ������������������������       �                     @        �       �                  S�2@z�G�z�?             @       �       �                   �<@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                 ���@���!pc�?             6@        ������������������������       �                      @        �       �                 �&B@z�G�z�?             4@       �       �                 ���@�q�q�?	             (@        ������������������������       �                      @        �       �                    �?���Q��?             $@       �       �                   �5@�q�q�?             "@        ������������������������       �                     �?        �       �                    9@      �?              @        ������������������������       �                     �?        ������������������������       �����X�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        �       �                   �0@�q�q�?+            �R@        �       �                    �?�����?             5@        ������������������������       �                      @        �       �                    �?�KM�]�?             3@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ��T?@�C��2(�?             &@       ������������������������       �                     @        �       �                    @z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ��l4@���3L�?             K@       �       �                 @3�@؀�:M�?            �B@        �       �                 ��}@r�q��?             (@        ������������������������       �                     @        �       �                    B@�<ݚ�?             "@       �       �                   �8@      �?              @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                 `f�%@�q�����?             9@       �       �                    4@�q�q�?             .@        ������������������������       �                     @        �       �                 ��l#@r�q��?             (@       �       �                    I@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                 @3�/@z�G�z�?             $@        ������������������������       �                     @        �       �                 pff0@���Q��?             @        �       �                    ;@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        
             1@        �       �                   �;@�%��5�?�            r@        �       �                    �?     ��?M             `@       �       �                    �?��E��?F            �\@       �       �                    @��z6��??             Y@        ������������������������       �                      @        �       �                    �?d}h���?>            �X@        �       �                    /@X�<ݚ�?             "@        ������������������������       �                      @        �       �                    �?և���X�?             @       �       �                    5@���Q��?             @        ������������������������       �                     �?        �       �                    8@      �?             @       �       �                 ���@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?NKF����?7            @V@       �       �                   �:@�P�����?1            �S@       �       �                    �?�?�'�@�?/             S@       �       �                   �2@4?,R��?,             R@        ������������������������       �                     &@        �       �                 0��A@��.��?&            �N@       �       �                   �5@(2��R�?%            �M@        �       �                    �?H�V�e��?             A@        ������������������������       �                     @        �       �                   �4@�������?             >@       �       �                   �3@R���Q�?             4@       �       �                 �?�@�θ�?             *@        ������������������������       �                     @        �       �                 `�8"@�q�q�?             "@        ������������������������       ����Q��?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                 ��L@���Q��?             $@        ������������������������       �                     @        ������������������������       �                     @        �       �                 ���@`2U0*��?             9@        �       �                 �&b@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     5@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?���Q��?             $@        ������������������������       �                     �?        �       �                 `f2@�q�q�?             "@       �       �                    +@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     ,@        ������������������������       �                     ,@        �       �                   �<@��	l�?f             d@       �       �                 ��) @XB���?:            �U@       ������������������������       �        '             M@        �       �                    �?ܷ��?��?             =@       �       �                 pf� @z�G�z�?
             .@        ������������������������       �                      @        �       �                 �T�C@$�q-�?	             *@       ������������������������       �                     $@        ������������������������       ��q�q�?             @        ������������������������       �        	             ,@        �                          �?�L���?,            �R@                                  ?@�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @                                 �?P�2E��?(            @P@                                 >@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@                                 �?h㱪��?$            �K@             	                  �E@ �q�q�?             H@       ������������������������       �                     >@        
                      P�@�����H�?             2@        ������������������������       �                      @                                �F@z�G�z�?             $@                              pf(@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �t�b��     h�h*h-K ��h/��R�(KMKK��h]�B        ~@      m@     �d@     �a@     �a@     �V@      O@     �M@      L@      C@      �?      2@      �?       @               @      �?                      0@     �K@      4@      $@      $@              @      $@      @       @      @      @      @      @              �?      @              @      �?              �?               @      @       @                      @     �F@      $@       @      @              �?       @       @       @                       @     �E@      @      >@      @      2@      @      2@      @       @              $@      @      @      @      @      @      @      @      @      �?       @      �?              �?       @              �?                       @      @                      �?      @                      @      (@              *@              @      5@      @      4@              &@      @      "@              "@      @              @      �?              �?      @              T@      @@      �?      ;@              3@      �?       @      �?       @      �?                       @              @     �S@      @      N@      @     �M@       @      7@              B@       @      1@       @       @              "@       @              �?      "@      �?      @               @      �?      �?      �?      �?              3@              �?      @              @      �?              3@              8@     �H@      1@      5@      �?      ,@      �?                      ,@      0@      @      0@      @      $@      @      @      �?      @              �?      �?      �?                      �?      @      @              @      @              @                      �?      @      <@      @      <@      �?      4@              @      �?      *@               @      �?      @              @      �?              @       @       @       @              @       @      �?              �?       @               @               @             �s@      W@     �L@      N@      @     �A@      @      :@      �?      $@              @      �?      @              @      �?      @      �?      @      �?                      @              �?      @      0@       @              @      0@      @       @               @      @      @      @      @      �?               @      @              �?       @      @      �?                       @              "@      I@      9@      3@       @       @              1@       @      @      �?              �?      @              $@      �?      @              @      �?              �?      @              ?@      7@      ,@      7@       @      $@              @       @      @      �?      @      �?      �?      �?                      �?              @      �?              (@      *@      $@      @              @      $@       @      @       @      @                       @      @               @       @              @       @      @       @      �?       @                      �?               @      1@             p@      @@     @Z@      7@     �V@      7@     @S@      7@               @     @S@      5@      @      @       @              @      @       @      @              �?       @       @       @      �?              �?       @                      �?      �?      �?      �?                      �?      R@      1@     �P@      *@     �P@      $@      O@      $@      &@             �I@      $@     �I@       @      ;@      @      @              7@      @      1@      @      $@      @      @              @      @       @      @      @              @              @      @              @      @              8@      �?      @      �?      @                      �?      5@                       @      @                      @      @      @              �?      @      @      �?      @              @      �?              @              ,@              ,@              c@      "@      U@      @      M@              :@      @      (@      @               @      (@      �?      $@               @      �?      ,@              Q@      @      @      @              @      @              O@      @      "@      �?              �?      "@             �J@       @      G@       @      >@              0@       @       @               @       @      �?       @               @      �?              @              @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�
HyhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B@F         |                   �'@4�<����?�           @�@               1                    �?��̇�?�             s@                                   �?Z��Yo��?+             O@                                   �?8�Z$���?             :@        ������������������������       �                     @                                  �2@��s����?             5@        ������������������������       �                     @               	                   �5@������?             1@        ������������������������       �                     �?        
                           9@     ��?
             0@        ������������������������       �                     �?                                   �?z�G�z�?	             .@                               ���@$�q-�?             *@        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                      @               0                    �?)O���?             B@              /                    �?�xGZ���?            �A@              .                    �?��.k���?             A@              '                   �=@��S���?             >@                                   @8�A�0��?             6@        ������������������������       �                     @                                   0@�����?             3@        ������������������������       �                     @               &                   �;@      �?             0@              #                 pf� @��
ц��?             *@              "                   �8@����X�?             @                               P��@���Q��?             @        ������������������������       �                      @                                   4@�q�q�?             @        ������������������������       �                     �?                !                 pff@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        $       %                    3@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        (       )                     @      �?              @        ������������������������       �                     @        *       +                    C@�q�q�?             @        ������������������������       �                     �?        ,       -                 `fV!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        2       G                    �?�C��2(�?�            @n@        3       F                 �y�#@�t����?#            �I@       4       =                  s�@ףp=
�?"             I@        5       <                   �7@�nkK�?             7@        6       ;                    �?؇���X�?             @       7       8                   �5@r�q��?             @        ������������������������       �                     @        9       :                 ���@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     0@        >       E                 ��(@PN��T'�?             ;@       ?       B                   �<@���y4F�?             3@       @       A                    �?�C��2(�?             &@       ������������������������       �ףp=
�?             $@        ������������������������       �                     �?        C       D                    >@      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        H       {                    �?�! �	��?x            �g@       I       z                    �?��Օ��?v            `g@       J       K                     @T�\�9�?u             g@        ������������������������       �                     :@        L       _                 �?�@ E�+0+�?e            �c@       M       ^                   @@@�ȉo(��?=            �V@       N       [                   �?@`Jj��?,             O@       O       P                   �7@P���Q�?*             N@        ������������������������       �                     <@        Q       R                 ���@     ��?             @@        ������������������������       �                      @        S       T                    ;@(;L]n�?             >@        ������������������������       �                     "@        U       Z                  sW@���N8�?             5@        V       Y                    =@�����H�?             "@       W       X                 pf�@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     (@        \       ]                   �@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     =@        `       y                    �?@�0�!��?(             Q@       a       f                 @3�@� y���?'            �P@        b       c                    :@�q�q�?             @        ������������������������       �                     �?        d       e                   �A@z�G�z�?             @        ������������������������       �                     @        ������������������������       �      �?              @        g       p                   �<@Xny��?"            �N@       h       k                   �3@��S�ۿ?            �F@        i       j                    2@"pc�
�?             &@       ������������������������       �                      @        ������������������������       ��q�q�?             @        l       m                 ��) @г�wY;�?             A@       ������������������������       �        
             4@        n       o                 pf� @@4և���?             ,@        ������������������������       �                     �?        ������������������������       �                     *@        q       x                 ��)"@      �?	             0@       r       w                   �@@$�q-�?             *@        s       v                 ��i @r�q��?             @       t       u                    ?@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        }                          @7i����?           �y@       ~                          @8��U��?�            @x@              �                    �?����?�            x@        �       �                     @<���D�?i            �d@       �       �                    �?�-.�1a�?J            �^@        ������������������������       �        %            �N@        �       �                     �?�g�y��?%             O@       �       �                    #@      �?             @@        ������������������������       �                      @        ������������������������       �                     >@        ������������������������       �                     >@        �       �                    @և���X�?             E@       �       �                 ��.@*O���?             B@        �       �                   �"@���|���?	             &@        ������������������������       �                      @        �       �                    �?�<ݚ�?             "@        ������������������������       �                     @        �       �                 ��*@���Q��?             @        ������������������������       �                     �?        �       �                 03�-@      �?             @        ������������������������       �                     �?        �       �                   �<@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 03�7@�+e�X�?             9@       �       �                   �=@�㙢�c�?             7@       �       �                    ;@      �?             0@        �       �                    �?      �?              @        �       �                    9@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?և���X�?             @       �       �                   �@@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   �>@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 ��D:@^(��I�?�            �k@       �       �                    @(N:!���?D            @Z@        �       �                     @؇���X�?             @       ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?��<D�m�?>            �X@        �       �                    �?�d�����?             3@       �       �                    �?@�0�!��?             1@       �       �                    =@$�q-�?             *@       �       �                    �?�����H�?	             "@       �       �                    �?r�q��?             @       �       �                 �R,@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                 �=/@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?�Fǌ��?0            �S@       �       �                   �*@�Ń��̧?             E@        �       �                 `fF)@�X�<ݺ?             2@        ������������������������       �                      @        �       �                   �;@      �?             0@       ������������������������       �                      @        �       �                    =@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     8@        ������������������������       �                    �B@        �                          �?
���n<�?C            �\@       �       �                 `f�B@h�|�`�?3            �U@        �       �                     �?�P�*�?             ?@       �       �                    �?����"�?             =@        �       �                 ��L@@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 `fF<@���Q��?             9@        �       �                    J@�eP*L��?             &@       �       �                 03k:@����X�?             @        ������������������������       �                      @        �       �                   @G@���Q��?             @       �       �                   @B@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   @>@����X�?             ,@        ������������������������       �                      @        �       �                   �J@�q�q�?             (@       �       �                   �>@z�G�z�?             $@        ������������������������       �                     @        �       �                   @B@���Q��?             @       �       �                   �@@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                 0�"K@�b��[��?            �K@        ������������������������       �                     &@        �       �                    �?~�4_�g�?             F@        �       �                    �?     ��?
             0@        �       �                   �8@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �H@�	j*D�?             *@       �       �                 �U�X@"pc�
�?             &@       �       �                 ���S@ףp=
�?             $@        ������������������������       �                     @        �       �                   �:@z�G�z�?             @        ������������������������       �                     @        �       �                 ��hU@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?����X�?             <@        ������������������������       �                     @        �       �                 `�jM@�q�q�?             8@        �       �                    ;@�q�q�?             (@        ������������������������       �                     �?        �       �                    >@�eP*L��?             &@       ������������������������       �      �?             $@        ������������������������       �                     �?                                   �?�8��8��?             (@                                �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @                              `fa@>���Rp�?             =@                               pA@�X����?             6@        ������������������������       �                     @                                 �?j���� �?
             1@       	      
                   +@�q�q�?	             .@        ������������������������       �                     @                               D�\@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @                                 �?ףp=
�?             4@        ������������������������       �                     @                                 @؇���X�?             ,@                              pf�C@���Q��?             @                                @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     "@        �t�bh�h*h-K ��h/��R�(KMKK��h]�B�        |@     �p@     `n@     �N@      7@     �C@      @      6@              @      @      1@              @      @      *@      �?              @      *@              �?      @      (@      �?      (@      �?                      (@       @              3@      1@      3@      0@      2@      0@      ,@      0@      *@      "@              @      *@      @      @              $@      @      @      @       @      @       @      @               @       @      �?      �?              �?      �?              �?      �?                       @      @      �?              �?      @              @              �?      @              @      �?       @              �?      �?      �?      �?                      �?      @              �?                      �?     �k@      6@     �F@      @     �F@      @      6@      �?      @      �?      @      �?      @              �?      �?              �?      �?              �?              0@              7@      @      .@      @      $@      �?      "@      �?      �?              @      @              @      @               @                      �?     �e@      0@     `e@      0@      e@      0@      :@             �a@      0@     �U@      @      M@      @     �L@      @      <@              =@      @               @      =@      �?      "@              4@      �?       @      �?      @      �?      @                      �?       @              (@              �?      �?              �?      �?              =@              L@      (@      L@      &@       @      @      �?              �?      @              @      �?      �?      K@      @      E@      @      "@       @       @              �?       @     �@@      �?      4@              *@      �?              �?      *@              (@      @      (@      �?      @      �?      @      �?      @                      �?       @              @                      @              �?       @              @             �i@     `i@     `g@      i@      g@      i@      4@      b@       @     @^@             �N@       @      N@       @      >@       @                      >@              >@      2@      8@      *@      7@      @      @               @      @       @      @              @       @              �?      @      �?      �?               @      �?       @                      �?      @      3@      @      3@      �?      .@      �?      @      �?       @               @      �?                      @               @      @      @      @      �?      @                      �?              @       @              @      �?      @                      �?     �d@      L@     @W@      (@      �?      @              @      �?      �?              �?      �?              W@      @      ,@      @      ,@      @      (@      �?       @      �?      @      �?      @      �?              �?      @               @              @              @               @       @       @                       @               @     �S@      �?     �D@      �?      1@      �?       @              .@      �?       @              @      �?              �?      @              8@             �B@             �Q@      F@     �H@     �B@      *@      2@      &@      2@      �?      @      �?                      @      $@      .@      @      @       @      @               @       @      @       @       @      �?       @      �?                      �?      @              @      $@               @      @       @       @       @              @       @      @      �?      @      �?                      @      �?               @               @              B@      3@      &@              9@      3@      @      &@      �?       @      �?                       @      @      "@       @      "@      �?      "@              @      �?      @              @      �?      �?      �?                      �?      �?               @              4@       @      @              0@       @      @      @              �?      @      @      @      @              �?      &@      �?      @      �?      @                      �?      @              6@      @      .@      @      @              $@      @      $@      @              @      $@      �?      $@                      �?               @      @              @              2@       @      @              (@       @      @       @      �?       @      �?                       @       @              "@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ���]hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B�D         <                    �?T�����?�           @�@                                ���=@ҳ�wY;�?O            �]@                                 �=@�^�����?)             O@                                  �?ڡR����?             �H@                                P�-@P���Q�?             4@        ������������������������       �                     &@               
                    �?�����H�?             "@               	                   �<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                ���@J�8���?             =@        ������������������������       �                     @                                @Q,@���Q��?             9@                               83##@��S���?	             .@                                  8@�z�G��?             $@        ������������������������       �                      @                                  �<@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @                                    �?z�G�z�?             $@                                �ܵ<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   �?      �?              @       ������������������������       �                     @                                �&2.@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        	             *@                ;                    �?�S����?&            �L@       !       "                    �?�2����?%            �K@       ������������������������       �                    �@@        #       $                 �EC@8�A�0��?             6@        ������������������������       �                     @        %       :                     �?�\��N��?             3@       &       3                    �?X�<ݚ�?             2@       '       2                   �D@�eP*L��?             &@       (       1                    �?�q�q�?             "@       )       .                    �?      �?              @       *       +                 ���Z@�q�q�?             @        ������������������������       �                      @        ,       -                 @�?t@      �?             @        ������������������������       �                      @        ������������������������       �                      @        /       0                 �̾w@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        4       5                 ��+T@և���X�?             @        ������������������������       �                     @        6       9                 �U�X@      �?             @        7       8                   �U@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        =       n                    �?bN�e�d�?v           ��@        >       E                     @������?m             e@        ?       @                    �?�"w����?6             S@       ������������������������       �        +            �N@        A       B                 ���`@��S�ۿ?             .@       ������������������������       �        	             (@        C       D                    8@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        F       c                    �?�û��|�?7             W@       G       N                 ��@D������?#            @P@        H       M                   �3@      �?	             0@        I       J                    1@���Q��?             @        ������������������������       �                     �?        K       L                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     &@        O       X                 Ь�#@ڡR����?            �H@       P       W                 @3�@\-��p�?             =@       Q       R                   �9@�<ݚ�?	             2@       ������������������������       �                     "@        S       T                    �?X�<ݚ�?             "@        ������������������������       �                      @        U       V                   �;@����X�?             @       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     &@        Y       \                    �?z�G�z�?             4@        Z       [                    4@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ]       ^                    �?r�q��?	             2@        ������������������������       �                     @        _       `                    ;@�θ�?             *@        ������������������������       �                      @        a       b                 03�1@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        d       m                    @�>����?             ;@       e       l                 @3�2@ףp=
�?             4@        f       k                    :@����X�?             @        g       h                   �#@�q�q�?             @        ������������������������       �                     �?        i       j                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             *@        ������������������������       �                     @        o       z                    !@�繠5�?	           �z@        p       q                     @П[;U��?             =@        ������������������������       �                     "@        r       s                     @��Q��?             4@        ������������������������       �                     @        t       u                    �?������?	             1@       ������������������������       �                     $@        v       y                    @և���X�?             @       w       x                    @z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        {                          �?�禺f��?�            �x@       |                         @S@dx@����?�            �u@       }       �                 ��$:@2Ǎ;�N�?�            �u@       ~       �                   �F@\�JЂ.�?�            `r@              �                  ��@���B��?�            pp@        �       �                     @ ,��-�?#            �M@        ������������������������       �        	             0@        �       �                 ��@�ʈD��?            �E@        �       �                    �?      �?              @        ������������������������       �                     @        �       �                 ���@z�G�z�?             @       �       �                    A@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �A@        �       �                   �<@��hJ,�?�            �i@       �       �                 �?$@8��8���?\             b@        �       �                 ��@���Q��?
             .@        �       �                    7@����X�?             @        ������������������������       �                      @        �       �                    �?���Q��?             @       ������������������������       �      �?             @        ������������������������       �                     �?        �       �                    6@      �?              @        ������������������������       �                      @        �       �                   �9@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                   �4@Du9iH��?R             `@        �       �                 pf� @"pc�
�?             6@        �       �                    �?���|���?             &@       �       �                   �3@�z�G��?             $@       �       �                 �?�@      �?              @        ������������������������       �                     @        �       �                   �1@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        	             &@        �       �                     @�f�¦ζ?B            �Z@        �       �                   �(@�C��2(�?             6@        ������������������������       �                     @        �       �                   �;@�r����?             .@       ������������������������       �        
             *@        ������������������������       �                      @        �       �                 м�5@@�)�n�?3            @U@       �       �                 ��) @F|/ߨ�?0            @T@       ������������������������       �                    �F@        �       �                 pf� @�X�<ݺ?             B@        ������������������������       �                     �?        �       �                    �?��?^�k�?            �A@        ������������������������       �                     @        �       �                    �?      �?             @@       �       �                 ���!@���N8�?             5@        �       �                    8@�q�q�?             @        ������������������������       �                     �?        �       �                   �;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             2@        ������������������������       �                     &@        �       �                 03�7@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 @3�@      �?+             N@        �       �                    �?���|���?             6@       �       �                    E@���Q��?             4@       �       �                   �?@�q�q�?             2@        �       �                    �?���Q��?             @        �       �                    >@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �>@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 �?�@�θ�?
             *@        ������������������������       �                     @        �       �                   �A@և���X�?             @       ������������������������       ����Q��?             @        ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                      @        �       �                     @>A�F<�?             C@       �       �                    �?�θ�?             :@       �       �                 `fF)@      �?
             0@        ������������������������       �                     @        �       �                   @B@���|���?             &@        �       �                    @@      �?             @        ������������������������       �                     �?        ������������������������       ����Q��?             @        �       �                   �3@z�G�z�?             @       ������������������������       �      �?             @        ������������������������       �                     �?        �       �                   �@@z�G�z�?             $@        �       �                   �>@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   �>@�8��8��?             (@        �       �                 ���"@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     ?@        �                            @r�z-��?"            �J@       �       �                   �;@f.i��n�?            �F@        �       �                    7@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                     �?      �?             D@       �       �                   �J@����>�?            �B@       �       �                   �>@J�8���?             =@        �       �                 `fF<@      �?              @       ������������������������       �                     @        �       �                   �<@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    D@؇���X�?             5@       �       �                   �B@�θ�?
             *@       �       �                    �?r�q��?	             (@       �       �                   �=@z�G�z�?             $@       �       �                 ��yC@�<ݚ�?             "@        �       �                   �A@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @                                 ;@      �?              @        ������������������������       �                     @                                 >@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @                                  @=QcG��?            �G@             	                   )@     ��?             @@        ������������������������       �                     �?        
                        �A@`Jj��?             ?@        ������������������������       �        	             .@                                 �?      �?	             0@        ������������������������       �                      @                                �B@؇���X�?             ,@                                 �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �                     .@        �t�bh�h*h-K ��h/��R�(KMKK��h]�B0       0|@     Pp@      E@     @S@     �@@      =@      4@      =@      �?      3@              &@      �?       @      �?       @      �?                       @              @      3@      $@      @              .@      $@      @       @      @      @               @      @      �?      @                      �?              @       @       @      �?      �?      �?                      �?      @      �?      @               @      �?       @                      �?      *@              "@      H@      "@      G@             �@@      "@      *@              @      "@      $@       @      $@      @      @      @      @      @      @       @      @               @       @       @       @                       @      �?      �?      �?                      �?              �?       @              @      @              @      @      �?      �?      �?      �?                      �?       @              �?                       @     �y@      g@     �L@     �[@      �?     �R@             �N@      �?      ,@              (@      �?       @               @      �?              L@      B@      ?@      A@       @      ,@       @      @              �?       @       @       @                       @              &@      =@      4@      9@      @      ,@      @      "@              @      @               @      @       @               @      @              &@              @      0@      �?      �?              �?      �?              @      .@              @      @      $@       @              �?      $@              $@      �?              9@       @      2@       @      @       @      �?       @              �?      �?      �?      �?                      �?      @              *@              @              v@     @R@      *@      0@              "@      *@      @              @      *@      @      $@              @      @      �?      @              @      �?               @             0u@     �L@     pr@      K@     pr@      J@     @p@      A@     �l@      A@     �K@      @      0@             �C@      @      @      @      @              �?      @      �?      �?              �?      �?                      @     �A@             �e@      >@      `@      .@      "@      @      @       @       @              @       @       @       @      �?              @      @       @               @      @              @       @              ^@      "@      2@      @      @      @      @      @      @      @      @              �?      @      �?                      @       @                      �?      &@             �Y@      @      4@       @      @              *@       @      *@                       @     �T@      @     �S@       @     �F@              A@       @              �?      A@      �?      @              ?@      �?      4@      �?       @      �?      �?              �?      �?              �?      �?              2@              &@              @      �?              �?      @             �F@      .@      ,@       @      (@       @      (@      @       @      @      �?      �?              �?      �?              �?       @      �?                       @      $@      @      @              @      @      @       @      �?      �?               @       @              ?@      @      4@      @      (@      @      @              @      @      @      @      �?               @      @      @      �?      @      �?      �?               @       @      �?       @      �?                       @      @              &@      �?       @      �?       @                      �?      "@              ?@             �A@      2@      ?@      ,@      �?      @      �?                      @      >@      $@      ;@      $@      3@      $@      �?      @              @      �?       @               @      �?              2@      @      $@      @      $@       @       @       @      @       @      @       @      @                       @      @              �?               @                      �?       @               @              @              @      @              @      @      �?      @                      �?               @      F@      @      =@      @              �?      =@       @      .@              ,@       @       @              (@       @       @       @       @                       @      $@              .@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�;hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM-huh*h-K ��h/��R�(KM-��h|�B@K         R                    �?�Qc�!�?�           @�@                                    @�<��S��?�            @o@                                  �?     �?Q             `@                                ��A@ 	��p�?             =@                                  @C@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     9@        	                        ���a@��:x�ٳ?@            �X@       
                           �?����ȫ�?7            �T@        ������������������������       �                    �C@                                   6@ qP��B�?            �E@                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                    �D@                                   !@@�0�!��?	             1@        ������������������������       �                     �?                                   �?      �?             0@       ������������������������       �                     *@                                   <@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?               O                 ���4@�p����?G            �^@                                 �1@�z��?8            @X@                                  �0@@4և���?             ,@       ������������������������       �                     $@                                �b&@      �?             @        ������������������������       �                     @        ������������������������       �                     �?               N                    @��q7L��?0            �T@               /                    �?L����?/            @T@        !       "                   �5@�eP*L��?             6@        ������������������������       �                     @        #       $                 ���@�q�q�?             2@        ������������������������       �                     @        %       &                    �?      �?	             (@        ������������������������       �                      @        '       .                 03�'@���Q��?             $@       (       -                 `f�@և���X�?             @       )       ,                    �?���Q��?             @       *       +                    9@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        0       M                    �?TV����?!            �M@       1       L                    @>4և���?             L@       2       K                    �?b�2�tk�?             K@       3       J                   @B@�E��
��?             J@       4       G                    �?(옄��?             G@       5       6                   �4@�G�z��?             D@        ������������������������       �                     @        7       @                 @3�@��
P��?            �A@        8       9                 ���@������?             .@        ������������������������       �                     @        :       =                 �&B@���|���?             &@        ;       <                   �7@      �?             @        ������������������������       �                     @        ������������������������       �                     @        >       ?                   �9@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        A       B                 `�X!@��Q��?             4@        ������������������������       �                     @        C       D                    ;@j���� �?	             1@       ������������������������       �                      @        E       F                 03�1@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        H       I                 03S1@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        P       Q                    �?`2U0*��?             9@        ������������������������       �                     �?        ������������������������       �                     8@        S       �                    �?��늓��?)           �|@       T       �                 ��$:@������?�             v@       U       n                    �?l���}��?�            pr@        V       m                 83�0@�t����?             A@       W       \                    9@���!pc�?            �@@        X       [                    �?r�q��?             @       Y       Z                 ��y@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ]       `                     @PN��T'�?             ;@        ^       _                 ���,@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        a       l                    ?@H%u��?             9@       b       k                 H�Z&@r�q��?
             2@       c       d                 ���@z�G�z�?	             .@        ������������������������       �                      @        e       j                   �<@�θ�?             *@       f       i                   @<@r�q��?             (@       g       h                   @@"pc�
�?             &@       ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        o       z                 ���@@�Žn��?�            Pp@        p       q                    �?�n`���?             ?@        ������������������������       �                     @        r       y                   �;@d}h���?             <@        s       t                 ��@�eP*L��?             &@        ������������������������       �                     @        u       v                    7@����X�?             @        ������������������������       �                     @        w       x                 �&b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        	             1@        {       �                    �?t��%�?�            �l@        |       �                   �=@`2U0*��?             9@       }       ~                   �:@P���Q�?
             4@        ������������������������       �                      @               �                 ��(@�X�<ݺ?	             2@       ������������������������       �$�q-�?             *@        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?������?�            �i@       �       �                     @8Fb����?~            @i@        �       �                   �;@(��+�?$            �N@        ������������������������       �                     8@        �       �                   �*@���@��?            �B@       �       �                 `f�)@l��
I��?             ;@        �       �                   @L@�����H�?             "@       ������������������������       �                     @        �       �                   �P@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    =@b�2�tk�?
             2@        ������������������������       �                     @        �       �                   �F@8�Z$���?	             *@       �       �                   @D@�<ݚ�?             "@       �       �                    @@      �?              @        ������������������������       �                      @        �       �                   @B@r�q��?             @       ������������������������       �z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        �       �                    �?�{"z;m�?Z            �a@       �       �                   �?@���}<S�?W            @a@       �       �                   �5@P���Q�??             Y@        �       �                 pf� @ �Cc}�?             <@       �       �                 �?$@r�q��?             2@        ������������������������       �                     @        �       �                   �4@���!pc�?             &@       �       �                 �?�@�����H�?             "@       ������������������������       �                     @        �       �                   �3@z�G�z�?             @       ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     $@        �       �                 pf� @������?-             R@       ������������������������       �        &             P@        �       �                   �8@      �?              @        ������������������������       �                     @        �       �                   �;@���Q��?             @        ������������������������       �                     �?        �       �                 ���"@      �?             @        ������������������������       �                     �?        �       �                   �<@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                 ��i @>A�F<�?             C@       �       �                   @@@R�}e�.�?             :@        �       �                 P�@���Q��?             $@        ������������������������       �                     @        �       �                 @3�@�q�q�?             @       ������������������������       �z�G�z�?             @        ������������������������       �                     �?        �       �                 �?�@      �?             0@       ������������������������       �                     $@        �       �                   �C@r�q��?             @        ������������������������       �                     @        �       �                   �G@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     (@        �       �                 @�$@�q�q�?             @        ������������������������       �                     �?        �       �                    9@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                     @TV����?,            �M@       �       �                    �?�"U����?'            �I@       �       �                   �>@r�qG�?$             H@        �       �                    �?r�q��?             8@        �       �                 ���<@�z�G��?             $@        ������������������������       �                     @        �       �                 ��>@      �?             @       �       �                   �E@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    K@����X�?             ,@       �       �                 `f�;@ףp=
�?             $@        ������������������������       �                     @        �       �                   `B@z�G�z�?             @        ������������������������       �                      @        �       �                   `H@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �Q@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 p�w@r�q��?             8@       �       �                   �;@�LQ�1	�?             7@        �       �                   �8@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?P���Q�?             4@        ������������������������       �                     @        �       �                    �?@4և���?             ,@       �       �                   �=@�C��2(�?	             &@       �       �                 `f�D@؇���X�?             @        �       �                   �A@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                 ��Ub@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                    ;@      �?              @        ������������������������       �                      @        �       �                    >@r�q��?             @        ������������������������       �      �?             @        ������������������������       �                      @        �                          �?�E��ӭ�?I             [@        �       �                 pVAH@�\��N��?             3@        �       �                 �&�)@�<ݚ�?             "@        �       �                 �x"@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   �5@z�G�z�?             $@        ������������������������       �                     �?                               p"�X@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?                                 �?�����L�?;            @V@                                �?��h!��?'            �L@        ������������������������       �                     @                                 +@�\�u��?#            �I@        ������������������������       �                      @                              03oY@&^�)b�?            �E@       	                      `fFJ@�p ��?            �D@       
                        �@@@4և���?             <@                                �?�����H�?             2@                               �>@8�Z$���?
             *@                                 @�8��8��?	             (@        ������������������������       �                      @                                �:@ףp=
�?             $@                             ��@z�G�z�?             @        ������������������������       �                      @                                �8@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@                                 C@�	j*D�?             *@                              `f�N@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @                                  �?      �?             @@        ������������������������       �                     @        !      ,                   @PN��T'�?             ;@       "      '                    @"pc�
�?             6@        #      &                   �?�q�q�?             @       $      %                  �B@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        (      )                   �?�KM�]�?
             3@       ������������������������       �                     .@        *      +                   @      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �t�b�@
     h�h*h-K ��h/��R�(KM-KK��h]�B�       �{@     �p@     �R@      f@      @     �^@       @      ;@       @       @               @       @                      9@      @     �W@      �?     @T@             �C@      �?      E@      �?      �?      �?                      �?             �D@      @      ,@      �?               @      ,@              *@       @      �?       @                      �?      Q@      K@      F@     �J@      �?      *@              $@      �?      @              @      �?             �E@      D@     �E@      C@      $@      (@      @              @      (@              @      @      @       @              @      @      @      @       @      @      �?      @              �?      �?       @      �?               @                      @     �@@      :@     �@@      7@     �@@      5@      ?@      5@      9@      5@      6@      2@      @              1@      2@      @      &@              @      @      @      @      @              @      @              �?      @      �?                      @      *@      @      @              $@      @       @               @      @              @       @              @      @      @                      @      @               @                       @              @               @      8@      �?              �?      8@              w@     �W@      r@      P@     p@      C@      8@      $@      8@      "@      �?      @      �?      @      �?                      @              �?      7@      @      �?      �?              �?      �?              6@      @      .@      @      (@      @       @              $@      @      $@       @      "@       @      @       @      @              �?                      �?      @              @                      �?      m@      <@      9@      @      @              6@      @      @      @              @      @       @      @              �?       @      �?                       @      1@              j@      6@      8@      �?      3@      �?       @              1@      �?      (@      �?      @              @              g@      5@     �f@      5@     �J@       @      8@              =@       @      3@       @       @      �?      @               @      �?              �?       @              &@      @              @      &@       @      @       @      @      �?       @              @      �?      @      �?      �?                      �?      @              $@              `@      *@     �_@      (@     �W@      @      9@      @      .@      @      @               @      @       @      �?      @              @      �?      �?      �?      @                       @      $@             �Q@       @      P@              @       @      @              @       @              �?      @      �?      �?               @      �?       @                      �?      ?@      @      3@      @      @      @              @      @       @      @      �?              �?      .@      �?      $@              @      �?      @               @      �?              �?       @              (@               @      �?      �?              �?      �?              �?      �?              @             �@@      :@      @@      3@      ?@      1@      &@      *@      @      @      @              @      @      @       @               @      @                      �?      @      $@      �?      "@              @      �?      @               @      �?       @      �?                       @      @      �?      @                      �?      4@      @      4@      @      �?       @      �?                       @      3@      �?      @              *@      �?      $@      �?      @      �?       @      �?       @                      �?      @              @              @                      �?      �?       @               @      �?              �?      @               @      �?      @      �?      @               @     �S@      >@      "@      $@      @       @      �?       @      �?                       @      @               @       @      �?              �?       @               @      �?             @Q@      4@     �D@      0@      @             �A@      0@               @     �A@       @     �A@      @      :@       @      0@       @      &@       @      &@      �?       @              "@      �?      @      �?       @               @      �?       @                      �?      @                      �?      @              $@              "@      @       @      @              @       @              @                       @      <@      @      @              7@      @      2@      @      �?       @      �?      �?      �?                      �?              �?      1@       @      .@               @       @               @       @              @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ� �thG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM1huh*h-K ��h/��R�(KM1��h|�B@L         p                     @�U��h��?�           @�@               #                    �?�(�k�I�?�             t@                                   �?���5��?1            �S@              	                    �?��Q��?             D@                                 �G@���N8�?             5@       ������������������������       �                     3@                                ,w�U@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        
                          �4@�����?             3@        ������������������������       �                      @                                �̾w@������?             1@                                  �?�r����?
             .@                                  A@8�Z$���?	             *@                                  �?�<ݚ�?             "@                               ���,@      �?              @        ������������������������       �                     �?                                   =@؇���X�?             @       ������������������������       �                     @                                `f `@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @                                   �?�˹�m��?             C@       ������������������������       �                     9@                                pVAH@�θ�?             *@        ������������������������       �                      @                                    �?�C��2(�?             &@       ������������������������       �                     @        !       "                   @K@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        $       %                    .@Υf���?�            �n@        ������������������������       �        
             *@        &       1                    �?J�����?�            �l@        '       (                    �?�d���?6            �U@       ������������������������       �        !             L@        )       0                   �;@`Jj��?             ?@        *       +                   �7@8�Z$���?	             *@        ������������������������       �                     �?        ,       -                   �8@�8��8��?             (@       ������������������������       �                     $@        .       /                 ���V@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     2@        2       o                    �?��a�2��?V             b@       3       j                    �?�ˡ�5��?U            �a@       4       5                   �:@HC>���?K            �^@        ������������������������       �                     3@        6       9                   �;@r�{o43�?=            �Y@        7       8                     �?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        :       i                 03�U@�����?:            �X@       ;       B                 `f�)@�"�q��?9            �W@        <       =                     �?���7�?             6@        ������������������������       �                     @        >       ?                   @L@      �?
             0@       ������������������������       �                     (@        @       A                   �P@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        C       h                   �J@��oh���?,            @R@       D       e                   �G@��6}��?%            �N@       E       T                     �?>���Rp�?"             M@       F       O                 �T!@@��R[s�?            �A@        G       N                    D@      �?             ,@       H       M                    @@X�<ݚ�?             "@       I       L                   @>@      �?              @       J       K                 `fF<@z�G�z�?             @       ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       ����Q��?             @        P       Q                   @K@�����?             5@       ������������������������       �                     *@        R       S                 03�M@      �?              @        ������������������������       �                      @        ������������������������       �                     @        U       d                   �E@��<b���?             7@       V       ]                   �*@�E��ӭ�?             2@        W       \                   @D@X�<ݚ�?             "@       X       Y                    @@r�q��?             @        ������������������������       �                     �?        Z       [                   @B@z�G�z�?             @       ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ^       _                   �7@�����H�?             "@        ������������������������       �                     @        `       c                   �:@r�q��?             @       a       b                   �@@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        f       g                     �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                     @        k       l                  x�F@P���Q�?
             4@       ������������������������       �                     .@        m       n                   �B@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        q       �                    �?؇>���?�            `x@        r       �                    �?@lܯ ��?N            �]@       s       �                    �?��z4���?,            @Q@        t       {                    �?     ��?             @@       u       x                    �?�LQ�1	�?             7@        v       w                   �+@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        y       z                 Ь* @�r����?	             .@       ������������������������       �                     *@        ������������������������       �                      @        |       �                 ���.@�q�q�?             "@        }       �                    �?      �?             @       ~                          �<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                 @3�2@4�B��?            �B@       �       �                 `�X!@      �?             @@       �       �                 ���@�<ݚ�?             2@        ������������������������       �                     �?        �       �                    ;@@�0�!��?             1@       �       �                 pf� @      �?             (@       �       �                   �9@�z�G��?             $@       �       �                   �6@      �?              @        �       �                    2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    7@և���X�?
             ,@       �       �                    �?      �?              @        �       �                  �#@z�G�z�?             @        ������������������������       �                      @        �       �                 �[$@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �#@�q�q�?             @        ������������������������       �                     �?        �       �                   �&@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?r�q��?             @       �       �                    A@z�G�z�?             @        ������������������������       �                      @        �       �                    I@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?`�Q��?"             I@        �       �                    �?և���X�?             @       �       �                 pF�-@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?^����?            �E@       �       �                 ��Y.@��H�}�?             9@        ������������������������       �                     "@        �       �                    �?     ��?             0@       �       �                    �?      �?             (@       �       �                 03�1@      �?              @       �       �                   �0@؇���X�?             @       �       �                    ;@      �?             @       �       �                 @3�/@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                 `fV6@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @r�q��?             2@        ������������������������       �                     @        �       �                    �?d}h���?
             ,@        ������������������������       �                     �?        �       �                   -@8�Z$���?	             *@        ������������������������       �                      @        ������������������������       �                     &@        �       0                  @@@vv@#_��?�            �p@       �       �                 �� @Xf1�
�?�            �l@        �       �                    6@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       #                   ?@�7�QJW�?�             l@       �                          @�����?�            �i@       �       �                    $@�r&��K�?{            `g@        ������������������������       �                     @        �       �                    �?D�N�dC�?w            �f@        �       �                    �?�J�4�?"             I@       �       �                    �?�*/�8V�?!            �G@       �       �                   �7@�C��2(�?             F@        �       �                    �?�<ݚ�?             "@       �       �                 xF*@����X�?             @       �       �                    5@      �?             @        �       �                 �{@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ���@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                 ���@ >�֕�?            �A@        ������������������������       �                     @        �       �                    �?@4և���?             <@       �       �                 ��(@�8��8��?             8@       �       �                 ���@�KM�]�?             3@        �       �                   @<@      �?              @       ������������������������       �z�G�z�?             @        ������������������������       �                     @        �       �                 03�@�C��2(�?             &@        ������������������������       �                      @        ������������������������       ������H�?             "@        ������������������������       �                     @        ������������������������       �                     @        �       �                   �1@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ��@�Ra����?U            �`@        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �                          �?�|K��2�?S             `@       �                         �:@`{��T��?D            @Y@       �       �                 ���@�.ߴ#�?)            �N@        �       �                 �&b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �                         �3@���#�İ?'            �M@        �       �                   �0@�C��2(�?             6@        �       �                 pFD!@      �?              @       �       �                 pf�@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �      �?             @        ������������������������       �                     @        �                          �2@@4և���?	             ,@        ������������������������       �                     @                              �?�@      �?              @       ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                    �B@                              ��) @R���Q�?             D@                             pb@؇���X�?             <@                              pf�@���Q��?             $@        ������������������������       �                     @        	      
                  �;@�q�q�?             @        ������������������������       �                      @        ������������������������       �      �?             @        ������������������������       �                     2@                              pf� @�q�q�?	             (@        ������������������������       �                      @                                �<@�z�G��?             $@                             �T�C@؇���X�?             @        ������������������������       �                     @        ������������������������       �      �?             @                              ���"@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                              pf� @h�����?             <@                                 �?ףp=
�?             $@                             P�@      �?              @        ������������������������       �                     @                                 8@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        
             2@                                  �?P���Q�?             4@       ������������������������       �                     ,@        !      "                pf�C@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        $      +                @3�@X�<ݚ�?	             2@       %      &                   �?���|���?             &@        ������������������������       �                     �?        '      (                  �@���Q��?             $@        ������������������������       �                     @        )      *                �?�@؇���X�?             @        ������������������������       �                     @        ������������������������       ��q�q�?             @        ,      -                ��i @؇���X�?             @        ������������������������       �                     @        .      /                d�6@@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �D@        �t�bh�h*h-K ��h/��R�(KM1KK��h]�B       �z@     �q@      a@      g@      1@     �N@      ,@      :@      �?      4@              3@      �?      �?      �?                      �?      *@      @               @      *@      @      *@       @      &@       @      @       @      @       @              �?      @      �?      @               @      �?              �?       @              �?              @               @                       @      @     �A@              9@      @      $@       @              �?      $@              @      �?      @      �?                      @      ^@      _@              *@      ^@     �[@       @     @U@              L@       @      =@       @      &@      �?              �?      &@              $@      �?      �?              �?      �?                      2@     �]@      :@     �]@      8@     �X@      7@      3@              T@      7@       @      @              @       @             �S@      4@     �S@      1@      5@      �?      @              .@      �?      (@              @      �?              �?      @             �L@      0@     �F@      0@      F@      ,@      :@      "@      @      @      @      @      @      @      @      �?      @      �?      �?                      @              �?      @       @      3@       @      *@              @       @               @      @              2@      @      *@      @      @      @      @      �?      �?              @      �?      @      �?      �?                      @       @      �?      @              @      �?      @      �?              �?      @              �?              @              �?       @               @      �?              (@                      @      3@      �?      .@              @      �?              �?      @                       @     `r@      X@     @P@      K@      ?@      C@      @      :@      @      4@      �?      @              @      �?               @      *@              *@       @              @      @      @      �?      �?      �?      �?                      �?       @                      @      9@      (@      4@      (@      ,@      @              �?      ,@      @      "@      @      @      @      @      �?      �?      �?      �?                      �?      @                       @       @              @              @       @      @      @      @      �?       @               @      �?              �?       @              �?       @              �?      �?      �?      �?                      �?      �?      @      �?      @               @      �?       @      �?                       @              �?      @              A@      0@      @      @      @       @      @                       @               @      ?@      (@      0@      "@      "@              @      "@      @      "@       @      @      �?      @      �?      @      �?      �?              �?      �?                       @              @      �?              �?      @              @      �?              @              .@      @      @              &@      @              �?      &@       @               @      &@             �l@      E@     �g@      E@       @      @       @                      @     @g@     �C@     @f@      =@     �c@      <@              @     �c@      7@      E@       @      E@      @      D@      @      @       @      @       @       @       @      �?      �?      �?                      �?      �?      �?              �?      �?              @               @             �@@       @      @              :@       @      6@       @      1@       @      @      �?      @      �?      @              $@      �?       @               @      �?      @              @               @      �?       @                      �?              @     @]@      .@      �?       @               @      �?              ]@      *@     @V@      (@      M@      @      �?      �?      �?                      �?     �L@       @      4@       @      @      �?      @      �?      �?              @      �?      @              *@      �?      @              @      �?      @              �?      �?     �B@              ?@      "@      8@      @      @      @      @               @      @               @       @       @      2@              @      @               @      @      @      @      �?      @              @      �?      �?       @      �?                       @      ;@      �?      "@      �?      @      �?      @              @      �?              �?      @               @              2@              3@      �?      ,@              @      �?              �?      @               @      $@      @      @      �?              @      @              @      @      �?      @               @      �?      �?      @              @      �?      @      �?                      @     �D@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ��1hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM	huh*h-K ��h/��R�(KM	��h|�B@B         d                     @r�����?�           @�@               7                  x#J@��J�fj�?�            �t@                                  (@n=�k��?�             l@        ������������������������       �        
             3@                                   @�ɭ�BR�?~            �i@        ������������������������       �                     "@                                   �?8�aW��?x            �h@               	                   �H@����e��?+            �P@       ������������������������       �        %             L@        
                           �?ףp=
�?             $@                                   �?�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?               *                     �?j��>��?M            ``@               )                 `f�B@θ	j*�?              J@                                ��>@��Zy�?            �C@                               ��$:@�	j*D�?             :@        ������������������������       �                     @                                   J@���|���?             6@                                 @@@և���X�?	             ,@                                   =@r�q��?             @                               �ܵ<@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @                                03k:@      �?              @        ������������������������       �                     @                                  @G@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        !       "                   @C@�	j*D�?	             *@        ������������������������       �                     @        #       $                   @H@և���X�?             @        ������������������������       �                      @        %       (                   @A@���Q��?             @       &       '                   �J@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     *@        +       6                    �?l{��b��?-            �S@       ,       -                 `f�)@��a�n`�?!             O@        ������������������������       �        
             1@        .       1                    =@�r����?            �F@        /       0                   �;@�E��ӭ�?	             2@       ������������������������       �                     *@        ������������������������       �                     @        2       3                   @D@ 7���B�?             ;@        ������������������������       �                     .@        4       5                    F@�8��8��?             (@        ������������������������       �      �?              @        ������������������������       �                     $@        ������������������������       �                     1@        8       c                    @����|e�?F             [@       9       :                    @�W;�E��?E            �Z@        ������������������������       �                     �?        ;       `                     �?�T`�[k�?D            �Z@       <       C                    �?Vβ���?@            @Y@       =       >                  "�b@��v$���?'            �N@       ������������������������       �                     H@        ?       B                    ;@$�q-�?	             *@        @       A                    8@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        D       Y                 `��`@      �?             D@       E       X                    �?���Q��?             >@       F       S                 ��hU@      �?             8@       G       N                    �?     ��?             0@        H       I                    �?      �?             @        ������������������������       �                      @        J       M                    �?      �?             @       K       L                 ��3Q@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        O       P                    8@z�G�z�?             $@        ������������������������       �                      @        Q       R                   @K@      �?              @        ������������������������       �                      @        ������������������������       �                     @        T       U                   �D@      �?              @        ������������������������       �                     @        V       W                   @G@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        Z       _                    �?z�G�z�?             $@       [       ^                    �?����X�?             @       \       ]                 @�?t@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        a       b                   PQ@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        e       �                    �?���皳�?�            �w@        f       �                    @�E1���?F            �Z@       g       �                   �=@�q�q�?E            @Z@       h                           �?�y�ʍ+�?=             W@        i       ~                 ��.@r٣����?            �@@       j       }                    �?�q�q�?             8@       k       |                 ���,@���!pc�?             6@       l       m                    �?z�G�z�?             4@        ������������������������       �                     @        n       {                    �?����X�?
             ,@       o       r                    4@�θ�?	             *@        p       q                   �0@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        s       z                 pF @"pc�
�?             &@       t       u                    9@ףp=
�?             $@        ������������������������       �                     �?        v       y                 �&B@�����H�?             "@       w       x                 ���@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     "@        �       �                 ���@�:�B��?'            �M@        ������������������������       �                     (@        �       �                   �<@��[�p�?!            �G@       �       �                    ;@:	��ʵ�?            �F@        �       �                    �?ҳ�wY;�?             1@       �       �                    +@�q�q�?             "@        ������������������������       �                      @        �       �                 ��&@և���X�?             @       �       �                    �?���Q��?             @       �       �                    5@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?@4և���?             <@        �       �                   @<@$�q-�?             *@       �       �                   @@�8��8��?             (@       ������������������������       �r�q��?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   `3@��S�ۿ?             .@       ������������������������       �                     &@        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     *@        ������������������������       �                      @        �       �                 03�1@��¤��?�             q@       �       �                 P��%@~X�<��?�             k@       �       �                    @ ��'^��?s            �g@       �       �                 @3�@��[�p�?r            �g@       �       �                 �?�@6�iL�?C            �]@       �       �                    �?�46<�?:             Y@       �       �                   �;@�����?8            �X@       �       �                 �1@�w��#��?             I@       �       �                    �?X�<ݚ�?             B@        ������������������������       �                     @        �       �                    7@8^s]e�?             =@       �       �                   �5@�X�<ݺ?
             2@       �       �                   �4@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        �       �                 ��@���!pc�?             &@        ������������������������       �                     @        �       �                    :@և���X�?             @       �       �                   �8@���Q��?             @       �       �                   �@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �@@4և���?	             ,@       �       �                 P�N@؇���X�?             @        ������������������������       �                      @        �       �                   �7@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   @@@      �?             H@       �       �                   �?@      �?             8@       ������������������������       �                     5@        ������������������������       �                     @        ������������������������       �                     8@        �       �                   �9@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?b�2�tk�?	             2@        ������������������������       �                     @        �       �                   �D@      �?             ,@       �       �                   �?@���|���?             &@        �       �                    :@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �A@      �?              @       ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �>@(N:!���?/            �Q@       �       �                    �?�X�<ݺ?$             K@       �       �                 @�!@ ��WV�?"             J@       �       �                    1@�7��?            �C@        ������������������������       �                     �?        �       �                   �;@P�Lt�<�?             C@        �       �                   �:@      �?             0@       ������������������������       �        
             .@        ������������������������       �                     �?        ������������������������       �                     6@        ������������������������       �                     *@        �       �                   �#@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?     ��?             0@        ������������������������       �                     @        �       �                    �?�8��8��?	             (@       �       �                 pf� @ףp=
�?             $@       �       �                   �@@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?�5��?             ;@        �       �                   �:@؇���X�?             ,@        �       �                    �?�q�q�?             @       �       �                 @3�/@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �*@�	j*D�?             *@        ������������������������       �                     @        �       �                   �/@ףp=
�?	             $@       ������������������������       �                     @        �       �                    (@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @4և����?$             L@        �       �                    @z�G�z�?             .@       �       �                 @3�4@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        �       �                 @3;:@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �                         �?@������?            �D@                                 �?��?^�k�?            �A@                                 �?�C��2(�?             &@                                ;@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     8@                                �A@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h*h-K ��h/��R�(KM	KK��h]�B�       �z@      r@      b@     �g@     �]@     �Z@              3@     �]@      V@      "@             @[@      V@      �?     @P@              L@      �?      "@      �?       @      �?                       @              �?      [@      7@     �A@      1@      6@      1@      2@       @      @              ,@       @      @       @      @      �?      @      �?      @                      �?       @              �?      @              @      �?      @      �?       @              �?       @              @      "@              @      @      @       @               @      @       @      �?              �?       @                       @      *@             @R@      @      L@      @      1@             �C@      @      *@      @      *@                      @      :@      �?      .@              &@      �?      �?      �?      $@              1@              :@     �T@      9@     �T@      �?              8@     �T@      5@      T@      �?      N@              H@      �?      (@      �?      @              @      �?                       @      4@      4@      (@      2@      (@      (@      &@      @      @      @       @              �?      @      �?      �?              �?      �?                       @       @       @       @              @       @               @      @              �?      @              @      �?      @      �?                      @              @       @       @      @       @       @       @       @                       @      @              @              @       @               @      @              �?             �q@     �X@     �Q@     �B@     �Q@     �A@     �L@     �A@       @      9@       @      0@      @      0@      @      0@              @      @      $@      @      $@      �?      �?              �?      �?               @      "@      �?      "@              �?      �?       @      �?       @              �?      �?      �?              @      �?              �?               @               @                      "@     �H@      $@      (@             �B@      $@     �B@       @      &@      @      @      @               @      @      @      @       @      �?       @               @      �?               @                       @       @              :@       @      (@      �?      &@      �?      @      �?      @              �?              ,@      �?      &@              @      �?      @                      �?               @      *@                       @     @j@      O@     �c@     �L@     �b@     �D@     �b@      D@     �U@      @@     �S@      5@     �S@      4@     �@@      1@      4@      0@              @      4@      "@      1@      �?      @      �?      @                      �?      $@              @       @              @      @      @      @       @       @       @               @       @              �?                       @      *@      �?      @      �?       @              @      �?      @                      �?      @             �F@      @      5@      @      5@                      @      8@              �?      �?              �?      �?              @      &@              @      @      @      @      @      �?       @      �?                       @      @       @      @       @       @                      @      O@       @     �I@      @      I@       @     �B@       @              �?     �B@      �?      .@      �?      .@                      �?      6@              *@              �?      �?              �?      �?              &@      @              @      &@      �?      "@      �?      @      �?              �?      @               @               @                      �?      &@      0@       @      (@       @      @       @       @               @       @                       @               @      "@      @              @      "@      �?      @              @      �?              �?      @             �I@      @      (@      @      "@      �?              �?      "@              @       @      @                       @     �C@       @      A@      �?      $@      �?      @      �?              �?      @              @              8@              @      �?              �?      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�JIhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B�A                            @������?�           @�@              ]                    �?����mA�?�           H�@                                    @V�a�� �?�             m@                                  �?P�2E��?S            @`@                                   �?`Jj��?;            @W@                                 �H@`2U0*��?             I@       ������������������������       �                    �C@                                �DD@"pc�
�?             &@        	       
                    K@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @                                  �;@�ʈD��?            �E@                                  �7@���|���?             &@                                   �?և���X�?             @        ������������������������       �                     �?                                   �?�q�q�?             @       ������������������������       �      �?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @@        ������������������������       �                    �B@               X                 ���4@j���� �??            �Y@              )                    �?:��?6            @V@                                0��@�I�w�"�?             C@        ������������������������       �                      @                                  �0@�z�G��?             >@        ������������������������       �                      @                                  �8@8�A�0��?             6@        ������������������������       �                     @               "                    �?������?
             1@                !                   �<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        #       (                    �?z�G�z�?             .@       $       '                    �?؇���X�?             ,@       %       &                  ��@z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        *       W                    �?j���� �?"            �I@       +       V                     @���H.�?!             I@       ,       9                   �5@և���X�?             �H@        -       8                    �?�z�G��?             $@       .       3                    0@�q�q�?             "@        /       0                    �?z�G�z�?             @        ������������������������       �                     @        1       2                   �&@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        4       5                 P��@      �?             @        ������������������������       �                     �?        6       7                 ��!@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        :       ;                   �@�99lMt�?            �C@        ������������������������       �                     @        <       M                 ��Y.@4���C�?            �@@       =       L                   �*@���Q��?             4@       >       K                    �?��.k���?             1@       ?       J                   P&@�n_Y�K�?	             *@       @       I                 ��l#@      �?             $@       A       B                 �?�@      �?              @        ������������������������       �                     �?        C       F                  SE"@����X�?             @       D       E                   �8@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        G       H                    I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        N       Q                    ;@8�Z$���?             *@        O       P                    9@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        R       S                 03�1@�C��2(�?             &@       ������������������������       �                     @        T       U                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        Y       \                 �A7@$�q-�?	             *@        Z       [                 `v�5@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        ^       �                    �?�v~y�/�?           |@       _       �                    �? ���	�?�            px@        `       m                   �;@�e�,��?%            �M@        a       l                 p"4W@      �?	             2@       b       c                      @�	j*D�?             *@        ������������������������       �                     @        d       e                 ��y@X�<ݚ�?             "@        ������������������������       �                     �?        f       g                   �0@      �?              @        ������������������������       �                      @        h       i                    8@r�q��?             @        ������������������������       �                     �?        j       k                 �0@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        n       �                 p�w@���?            �D@       o       �                   �G@R���Q�?             D@       p       �                   �=@��hJ,�?             A@       q       ~                   �<@�+$�jP�?             ;@       r       }                 03SA@      �?             8@       s       |                   @<@     ��?             0@       t       {                    �?z�G�z�?             .@       u       v                      @d}h���?             ,@        ������������������������       �                     �?        w       x                 ���@8�Z$���?
             *@        ������������������������       �                     @        y       z                   @@z�G�z�?             $@       ������������������������       �����X�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @               �                 ���1@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �H@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 �TL@��x���?�            �t@       �       �                     �?���1���?�            �s@        �       �                   @J@���y4F�?             C@       �       �                   `G@      �?             @@       �       �                 ��yC@�>4և��?             <@       �       �                   �<@�E��ӭ�?             2@        �       �                   `@@և���X�?             @       ������������������������       �                     @        �       �                   �A@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �B@�C��2(�?             &@        �       �                    @@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        �       �                   �H@      �?             @        ������������������������       �                      @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �:@��ׄ��?�            `q@        �       �                     @hl �&�?=             W@        ������������������������       �                     0@        �       �                   �0@p�|�i�?2             S@        �       �                 pf�@�q�q�?             @        ������������������������       �                     �?        �       �                 pFD!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 @33@��pBI�?/            @R@        ������������������������       �                     �?        �       �                    �?�k~X��?.             R@       �       �                 ���@ �.�?Ƞ?'             N@        �       �                    6@z�G�z�?             @        ������������������������       �                      @        �       �                 �&b@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        #            �K@        ������������������������       �                     (@        �       �                   �;@�I�,ѽ�?o            @g@        �       �                 ���%@      �?             $@        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?h�V���?k             f@       �       �                     @���(`�?j            �e@        �       �                   @N@P���Q�?             D@       �       �                    �?P�Lt�<�?             C@        ������������������������       �                     �?        �       �                   �4@�?�|�?            �B@       ������������������������       �                     8@        �       �                    �?$�q-�?             *@        ������������������������       �                     @        �       �                   �@@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?pH����?P            �`@       �       �                   �C@�����H�?K            �_@       �       �                    �?L紂P�?;            �Y@        �       �                   �<@�����?             5@       ������������������������       �        
             1@        �       �                    >@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                 �?�@PN��T'�?.            @T@        �       �                    =@`Jj��?             ?@       �       �                  sW@      �?
             0@        �       �                 pf�@�q�q�?             @        ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                     $@        ������������������������       �                     .@        �       �                   �<@z�G�z�?             I@       �       �                 pf� @ףp=
�?             >@       �       �                 ��) @z�G�z�?	             .@       ������������������������       �                     (@        ������������������������       �                     @        ������������������������       �                     .@        �       �                   @@@��Q��?             4@       �       �                 @3�@�eP*L��?             &@        ������������������������       �                      @        �       �                 ���"@�q�q�?             "@       �       �                 ��i @؇���X�?             @       �       �                    ?@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                 @3�@�<ݚ�?             "@        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     8@        ������������������������       �                      @        ������������������������       �                      @        �       �                    9@     ��?
             0@        ������������������������       �                      @        �       �                   �C@X�Cc�?             ,@       �       �                     @�	j*D�?             *@        ������������������������       �                      @        �       �                    >@"pc�
�?             &@       �       �                    ;@���Q��?             @        ������������������������       �                     �?        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    (@�BbΊ�?&             M@        ������������������������       �        
             *@        �                       @�:x@`Ӹ����?            �F@       �       �                    �?`���i��?             F@       ������������������������       �                     >@        �       �                    @@@4և���?             ,@        ������������������������       �                      @        �       �                    �?r�q��?             @        ������������������������       �                     �?        �                         �g@z�G�z�?             @                                  �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?                              hf�2@�g�y��?             ?@        ������������������������       �                     �?        ������������������������       �                     >@        �t�b��	     h�h*h-K ��h/��R�(KMKK��h]�Bp        |@     `p@     @z@     Pp@      H@      g@      @      _@      @     �U@       @      H@             �C@       @      "@       @      �?       @                      �?               @      @     �C@      @      @      @      @              �?      @       @       @       @       @                      @              @@             �B@      E@      N@      >@     �M@      "@      =@               @      "@      5@               @      "@      *@      @              @      *@      �?      �?      �?                      �?      @      (@       @      (@       @       @       @                       @              @      �?              5@      >@      5@      =@      5@      <@      @      @      @      @      @      �?      @              �?      �?      �?                      �?       @       @              �?       @      �?       @                      �?      �?              ,@      9@              @      ,@      3@      (@       @      "@       @      @       @      @      @      @      @      �?               @      @      �?      @      �?                      @      �?      �?      �?                      �?       @                      @      @              @               @      &@      �?      �?              �?      �?              �?      $@              @      �?      @      �?                      @              �?              �?      (@      �?      @      �?      @                      �?      "@             @w@     @S@     �t@      O@      D@      3@      "@      "@      @      "@              @      @      @      �?              @      @       @              �?      @              �?      �?      @      �?                      @      @              ?@      $@      ?@      "@      =@      @      6@      @      5@      @      *@      @      (@      @      &@      @              �?      &@       @      @               @       @      @       @      @              �?              �?               @              �?       @               @      �?              @               @      @              @       @                      �?     r@     �E@     �q@      A@      >@       @      8@       @      7@      @      *@      @      @      @              @      @      �?      @                      �?      $@      �?      @      �?      @                      �?      @              $@              �?      @               @      �?      �?              �?      �?              @             �o@      :@     @V@      @      0@             @R@      @       @      �?      �?              �?      �?              �?      �?             �Q@       @              �?     �Q@      �?     �M@      �?      @      �?       @               @      �?       @                      �?     �K@              (@             `d@      7@      @      @              @      @             �c@      2@     �c@      0@      C@       @     �B@      �?      �?              B@      �?      8@              (@      �?      @              @      �?              �?      @              �?      �?              �?      �?              ^@      ,@      \@      ,@      V@      ,@      3@       @      1@               @       @               @       @             @Q@      (@      =@       @      ,@       @      @       @      @              �?       @      $@              .@              D@      $@      ;@      @      (@      @      (@                      @      .@              *@      @      @      @               @      @      @      @      �?      @      �?      @                      �?      @                       @      @       @       @       @      @              8@               @                       @      @      "@       @              @      "@      @      "@       @               @      "@       @      @              �?       @       @              @      �?             �E@      .@              *@     �E@       @     �E@      �?      >@              *@      �?       @              @      �?      �?              @      �?      �?      �?              �?      �?              @                      �?      >@      �?              �?      >@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ��NhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B@D         j                     @Dl���v�?�           @�@               '                 ���<@r�q��?�             u@                                  @p�
�+�?g            �e@        ������������������������       �                     $@               "                    �?��P��?`            �d@                                  �?���f��?K            �_@                                   �?�}�+r��?             C@       ������������������������       �                     ?@        	       
                    �?����X�?             @        ������������������������       �                     �?                                  �7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @               !                    �?`���i��?2             V@                               ��$:@���Hx�?*             R@                                  &@�1�`jg�?            �K@                                  �7@���!pc�?             &@                                  �1@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     F@                                   �?������?             1@        ������������������������       �                     @                                   �J@����X�?
             ,@                                 @G@X�<ݚ�?             "@                               03k:@����X�?             @        ������������������������       �                     �?                                  @B@r�q��?             @        ������������������������       �                     �?        ������������������������       �z�G�z�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     0@        #       $                    �?���y4F�?             C@       ������������������������       �                     9@        %       &                    1@�n_Y�K�?             *@        ������������������������       �                     @        ������������������������       �                      @        (       W                 03?U@��4�-�?e            @d@       )       6                   �;@x�K��?B            �Y@        *       +                    2@�+$�jP�?             ;@        ������������������������       �                     "@        ,       3                     �?�E��ӭ�?             2@       -       2                 Ј@S@؇���X�?
             ,@       .       /                    �?$�q-�?	             *@       ������������������������       �                     "@        0       1                   �4@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        4       5                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        7       8                    �?��S���?0            �R@        ������������������������       �                     =@        9       F                    �?�5��
J�?             G@        :       ?                   �G@      �?
             0@       ;       >                   �A@���!pc�?             &@        <       =                    @@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        @       E                    �?���Q��?             @       A       B                   �J@�q�q�?             @        ������������������������       �                     �?        C       D                   �L@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        G       R                    �?r�q��?             >@       H       Q                     �?"pc�
�?             6@       I       P                 ��yC@��s����?             5@        J       O                   �<@      �?              @       K       L                   `@@z�G�z�?             @        ������������������������       �                      @        M       N                   �A@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        	             *@        ������������������������       �                     �?        S       V                  x�N@      �?              @        T       U                   @@@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        X       i                    @d��0u��?#             N@       Y       Z                     @&y�X���?"             M@        ������������������������       �                     @        [       d                    �?H�ՠ&��?!             K@       \       ]                    �?�n`���?             ?@       ������������������������       �                     5@        ^       _                   �7@���Q��?             $@        ������������������������       �                     @        `       a                 Ј�V@և���X�?             @        ������������������������       �                      @        b       c                   @E@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        e       f                    @�nkK�?             7@       ������������������������       �        
             4@        g       h                    5@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        k                        ��Y7@�*/�8V�?�            �w@       l       �                    �?Y!8�D�?�            �s@        m       �                    �?�ģ�a@�?:            @U@       n                          �5@�O�y���?2            �R@        o       ~                    �?�X����?             6@       p       {                    �?j���� �?             1@       q       t                    �?���Q��?
             .@        r       s                    0@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        u       x                    3@X�<ݚ�?             "@       v       w                    0@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        y       z                   �4@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        |       }                    %@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @H(���o�?#            �J@        �       �                   �9@��2(&�?             6@        �       �                 ��@�z�G��?             $@        ������������������������       �                     @        �       �                   �6@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        	             (@        �       �                    3@�g�y��?             ?@       �       �                    �?և���X�?             <@        ������������������������       �                     �?        �       �                   �:@X�<ݚ�?             ;@        ������������������������       �                     @        �       �                 ��1@�eP*L��?             6@       �       �                    �?�q�q�?             2@       �       �                    �?d}h���?             ,@        �       �                    =@�q�q�?             @        ������������������������       �                     �?        �       �                   �>@z�G�z�?             @        �       �                 @3#%@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                   @B@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?z�G�z�?             $@        �       �                 ���.@���Q��?             @        �       �                   �<@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    +@d{���2�?�            @m@        ������������������������       �                      @        �       �                    �?&^�r���?�            @l@       �       �                    �?�uX��?�             k@        �       �                    �?¦	^_�?             ?@       �       �                 �� @�+e�X�?             9@       �       �                 ��y@��+7��?             7@        ������������������������       �                     �?        �       �                    9@���!pc�?             6@        ������������������������       �                      @        �       �                 ���@z�G�z�?             4@        ������������������������       �                     @        �       �                   �=@������?
             1@       �       �                   �<@�	j*D�?             *@       �       �                   @<@"pc�
�?             &@       �       �                   @@�<ݚ�?             "@       ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                 ��&@      �?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �>@��� ��?{            @g@       �       �                    �?DS���|�?Z             a@        �       �                  s�@�����?             5@        ������������������������       �                     @        �       �                    �?�r����?             .@       ������������������������       �"pc�
�?             &@        ������������������������       �                     @        �       �                    �?ܷ��?��?O             ]@       �       �                    �?hdpZ�L�?L            @\@       �       �                   �;@�KM�]�?A            �W@       �       �                 ��@@�r-��?(            �M@        ������������������������       �                      @        �       �                 ��L@���5��?'            �L@        �       �                    4@���!pc�?             6@        ������������������������       �                      @        �       �                   �5@և���X�?
             ,@        �       �                  s@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �&b@�<ݚ�?             "@        ������������������������       �                      @        �       �                 03S@����X�?             @        ������������������������       �                     �?        �       �                 �?$@r�q��?             @        ������������������������       �                      @        �       �                   �9@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 ��Y @��?^�k�?            �A@       �       �                   �1@      �?             0@        ������������������������       �      �?              @        ������������������������       �                     ,@        ������������������������       �                     3@        �       �                 ��) @������?             B@       ������������������������       �                     ;@        �       �                 pf� @�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        �       �                 pf�'@�����H�?             2@        �       �                 ��@      �?              @        ������������������������       �                     @        �       �                   �9@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     @        �       �                    �?�����?!            �H@       �       �                    �?��<b���?             G@       �       �                   @@@>��C��?            �E@        �       �                   �?@�eP*L��?             &@        ������������������������       �                     �?        �       �                 @3�@      �?             $@       �       �                 �?�@      �?              @        ������������������������       �                     �?        ������������������������       �և���X�?             @        ������������������������       �                      @        �       �                 �?�@      �?             @@       ������������������������       �                     4@        �       �                 @3�@�q�q�?             (@        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                  �v6@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @                                 �?l�b�G��?'            �L@        ������������������������       �                     5@                                 �?�����H�?             B@        ������������������������       �                     @                                 �?      �?             @@                                �A@և���X�?             @             
                   �?���Q��?             @             	                   >@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @                                 @`2U0*��?             9@                                 @z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     4@        �t�bh�h*h-K ��h/��R�(KMKK��h]�B        {@     `q@     @c@     �f@     @Y@     @R@      $@             �V@     @R@     �T@     �E@       @      B@              ?@       @      @              �?       @      @       @                      @     @T@      @     @P@      @      J@      @       @      @       @      @       @                      @      @              F@              *@      @      @              $@      @      @      @      @       @              �?      @      �?      �?              @      �?               @      @              0@               @      >@              9@       @      @              @       @             �J@     @[@      D@      O@      @      6@              "@      @      *@       @      (@      �?      (@              "@      �?      @      �?                      @      �?              @      �?              �?      @             �A@      D@              =@     �A@      &@      $@      @       @      @      �?      @              @      �?              @               @      @       @      �?      �?              �?      �?              �?      �?                       @      9@      @      2@      @      1@      @      @      @      �?      @               @      �?       @      �?                       @      @              *@              �?              @      �?       @      �?       @                      �?      @              *@     �G@      &@     �G@      @              @     �G@      @      9@              5@      @      @      @              @      @       @              �?      @              @      �?              �?      6@              4@      �?       @      �?                       @       @             �q@      X@     `l@      W@      B@     �H@      A@     �D@      .@      @      $@      @      "@      @      @      �?              �?      @              @      @      �?      @      �?                      @      @      �?      @                      �?      �?      �?              �?      �?              @              3@      A@      @      3@      @      @              @      @      @              @      @                      (@      0@      .@      0@      (@      �?              .@      (@      @              $@      (@      @      (@      @      &@       @      @      �?              �?      @      �?       @      �?                       @               @      �?      @              @      �?              @      �?              �?      @              @                      @       @       @       @      @       @      �?       @                      �?               @              @     �g@     �E@               @     �g@     �A@      g@     �@@      6@      "@      3@      @      1@      @      �?              0@      @               @      0@      @      @              *@      @      "@      @      "@       @      @       @      @       @      @               @                       @      @               @              @      @      @                      @     @d@      8@     �^@      ,@      3@       @      @              *@       @      "@       @      @              Z@      (@     @Y@      (@     @U@      $@      I@      "@               @      I@      @      0@      @       @               @      @      �?      @      �?                      @      @       @       @              @       @              �?      @      �?       @              @      �?      @                      �?      A@      �?      .@      �?      �?      �?      ,@              3@             �A@      �?      ;@               @      �?              �?       @              0@       @      @       @      @              �?       @               @      �?              $@              @             �C@      $@      B@      $@     �@@      $@      @      @              �?      @      @      @      @      �?              @      @               @      <@      @      4@               @      @              @       @              @              @              @       @      @                       @     �J@      @      5@              @@      @      @              <@      @      @      @       @      @      �?      @      �?       @              �?      �?               @              8@      �?      @      �?      @                      �?      4@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ2�3hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM'huh*h-K ��h/��R�(KM'��h|�B�I         �                  x#J@l��n�?�           @�@              U                    �?��*?L�?o           `�@               T                    @z�t���?o             h@                                   @V���#�?l            �g@                                  �H@P�2E��?&            @P@                                 �8@ _�@�Y�?"             M@                                   �? 7���B�?             ;@              	                   �7@@4և���?	             ,@       ������������������������       �                     "@        
                            �?z�G�z�?             @        ������������������������       �                      @                                  �3@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     *@        ������������������������       �                     ?@                                  �I@����X�?             @                                03�3@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @               /                    �?l��TO��?F            @_@               .                 �?�-@�E��ӭ�?             K@              -                    �?��]�T��?            �D@                                 �5@�����?             C@                                   0@      �?             $@                                P��+@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @               ,                    �?      �?             <@               !                    �?�<ݚ�?             ;@        ������������������������       �                     @        "       #                    9@��+7��?             7@        ������������������������       �                      @        $       %                 ���@����X�?             5@        ������������������������       �                     @        &       +                 pF @�t����?             1@       '       (                 ���@      �?
             0@        ������������������������       �                     @        )       *                 �&B@$�q-�?             *@       ������������������������       �ףp=
�?             $@        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     *@        0       Q                    �?.}Z*�?'            �Q@       1       P                 �̼6@և���X�?             L@       2       O                    �?�eP*L��?             F@       3       4                 ���@����e��?            �@@        ������������������������       �                     @        5       D                    �?�q�q�?             >@       6       C                 ��l#@z�G�z�?             4@       7       8                 �&B@      �?             0@        ������������������������       �                      @        9       <                 P�@����X�?
             ,@        :       ;                    4@      �?             @        ������������������������       �                      @        ������������������������       �                      @        =       B                    I@z�G�z�?             $@       >       ?                    9@�����H�?             "@        ������������������������       �                     @        @       A                 @3�@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        E       H                    9@���Q��?             $@        F       G                    6@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        I       N                   �@@���Q��?             @       J       M                   �=@      �?             @       K       L                    ;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     (@        R       S                 ���)@z�G�z�?             .@        ������������������������       �                     @        ������������������������       �                     (@        ������������������������       �                     @        V       Y                    $@ m��R��?            �x@        W       X                    @D�n�3�?             3@       ������������������������       �        	             &@        ������������������������       �                      @        Z       y                     �?PcG���?�            �w@        [       \                   �;@6�iL�?!            �M@        ������������������������       �                      @        ]       ^                 ��$:@P̏����?             �L@        ������������������������       �                     "@        _       x                    �?�q�q�?             H@       `       a                 03k:@�X����?             F@        ������������������������       �                     @        b       q                 �TaA@���� �?            �D@       c       p                   �>@     ��?             @@       d       k                    �?�q�q�?             8@        e       f                 �ܵ<@      �?              @        ������������������������       �                     @        g       j                    �?      �?             @       h       i                   �E@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        l       m                   �<@      �?	             0@        ������������������������       �                     @        n       o                   �Q@r�q��?             (@       ������������������������       �                     $@        ������������������������       �                      @        ������������������������       �                      @        r       s                    �?X�<ݚ�?             "@        ������������������������       �                     @        t       w                   @B@r�q��?             @       u       v                 `f�D@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        z       �                    &@��3֞�?�            �s@       {       �                   �0@�F�1G�?�            �j@        |       �                    �?���Q��?             $@       }       �                 pFD!@      �?              @        ~                        pf�@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                   @N@L紂P�?            �i@       �       �                    �?0w-!��?}             i@       �       �                    �? ���3�?{            �h@        �       �                 ���@��2(&�?             F@        ������������������������       �                     $@        �       �                    �?@�0�!��?             A@       �       �                   @@z�G�z�?             4@       �       �                    5@�θ�?             *@        ������������������������       �                     @        ������������������������       �                     $@        �       �                    @@؇���X�?             @       �       �                   �<@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?؇���X�?	             ,@       �       �                   �=@8�Z$���?             *@       �       �                  s�@����X�?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?��}���?b            @c@       �       �                   �:@8F�V�?]            `b@        �       �                   �4@`'�J�?#            �I@        ������������������������       �                     2@        �       �                     @�FVQ&�?            �@@        ������������������������       �                     �?        �       �                 �1@      �?             @@        �       �                   �5@8�Z$���?	             *@        �       �                  s@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ���@�C��2(�?             &@        �       �                   �8@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     3@        �       �                   �;@     ��?:             X@        ������������������������       �                     @        �       �                   @@@*
;&���?7             W@       �       �                   �>@d}h���?              L@       �       �                   �<@�*/�8V�?            �G@       �       �                     @$�q-�?            �C@        ������������������������       �                     �?        �       �                 ��) @�˹�m��?             C@       �       �                  sW@�X�<ݺ?             B@        �       �                 pf�@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �      �?             @        ������������������������       �                     ;@        �       �                 �̜!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �=@      �?              @        �       �                 �̌!@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   �?@�<ݚ�?             "@        ������������������������       �                     @        �       �                 ��I @�q�q�?             @       �       �                 �?�@z�G�z�?             @       �       �                   �@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                     @�X�<ݺ?             B@        ������������������������       �                     @        �       �                   �E@      �?             @@       ������������������������       �                     3@        �       �                   �F@8�Z$���?	             *@        �       �                 @3�@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     @        ������������������������       �                      @        �       �                     @      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?b �57�?I            �Y@        �       �                    =@d}h���?             <@       �       �                    �?����X�?             5@       �       �                    �?     ��?             0@       �       �                     @���!pc�?             &@        �       �                 `��,@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                 ��$1@؇���X�?             @        ������������������������       �                     @        �       �                    �?�q�q�?             @       �       �                   �2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                  �v6@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    ?@�}��L�?6            �R@        ������������������������       �                    �B@        �       �                 039@P�Lt�<�?             C@       ������������������������       �                     :@        �       �                    �?�8��8��?	             (@       �       �                    �?؇���X�?             @        ������������������������       �                     @        �       �                   �@@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       $                    @x�����?M             _@       �                       ��LY@��h!��?D            �\@       �                         �P@d�;lr�?'            �O@       �       �                    �?f>�cQ�?&            �N@       ������������������������       �                    �D@        �       �                    �?�G�z��?             4@        ������������������������       �                      @        �                          �?b�2�tk�?             2@       �       �                   �;@     ��?             0@        ������������������������       �                     @        �                          �?�q�q�?
             (@                                  �?      �?             @                             ���S@�q�q�?             @        ������������������������       �                     �?                                @C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?                                 �?      �?              @                                E@և���X�?             @       	      
                `f�N@      �?             @        ������������������������       �                      @                              03�S@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @                                 �?j���� �?            �I@                             03c@z�G�z�?             >@                              ���a@      �?             0@       ������������������������       �                     "@                                �7@؇���X�?             @                                (@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             ,@              !                   �?����X�?             5@                                 �?d}h���?             ,@                               �?@      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        "      #                  �d@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        %      &                   �?�z�G��?	             $@        ������������������������       �                     @        ������������������������       �                     @        �t�bh�h*h-K ��h/��R�(KM'KK��h]�Bp       {@     pq@     �x@     @h@     @P@      `@      O@      `@      @      O@      �?     �L@      �?      :@      �?      *@              "@      �?      @               @      �?       @      �?                       @              *@              ?@       @      @       @      �?              �?       @                      @     �M@     �P@      .@     �C@      .@      :@      (@      :@      @      @      �?      @              @      �?              @              @      5@      @      5@              @      @      1@               @      @      .@      @               @      .@      �?      .@              @      �?      (@      �?      "@              @      �?              �?              @                      *@      F@      ;@      @@      8@      4@      8@      4@      *@              @      4@      $@      0@      @      (@      @       @              $@      @       @       @       @                       @       @       @       @      �?      @              @      �?              �?      @                      �?      @              @      @      �?      @      �?                      @      @       @      @      �?      �?      �?      �?                      �?       @                      �?              &@      (@              (@      @              @      (@              @             �t@     �P@       @      &@              &@       @             t@     �K@     �E@      0@               @     �E@      ,@      "@              A@      ,@      >@      ,@              @      >@      &@      9@      @      1@      @      @      �?      @              @      �?      �?      �?              �?      �?               @              $@      @              @      $@       @      $@                       @       @              @      @              @      @      �?       @      �?              �?       @              @              @             `q@     �C@     �f@      @@      @      @      @      @      �?      @      �?                      @      @               @              f@      <@     �e@      :@     �e@      :@      C@      @      $@              <@      @      0@      @      $@      @              @      $@              @      �?       @      �?       @                      �?      @              (@       @      &@       @      @       @      �?              @       @      @              �?             �`@      4@     �_@      4@     �H@       @      2@              ?@       @      �?              >@       @      &@       @      �?      �?      �?                      �?      $@      �?      @      �?              �?      @              @              3@             �S@      2@              @     �S@      ,@      F@      (@      E@      @      B@      @      �?             �A@      @      A@       @      @       @      @               @       @      ;@              �?      �?              �?      �?              @       @      �?       @      �?                       @      @               @      @              @       @      @      �?      @      �?      �?              �?      �?                      @      �?              A@       @      @              >@       @      3@              &@       @       @       @               @       @              "@              @               @               @       @               @       @              X@      @      6@      @      .@      @      *@      @       @      @       @       @               @       @              @      �?      @               @      �?      �?      �?      �?                      �?      �?              @               @      @       @                      @      @             �R@      �?     �B@             �B@      �?      :@              &@      �?      @      �?      @               @      �?              �?       @              @             �C@     @U@      @@     �T@      &@      J@      "@      J@             �D@      "@      &@       @              @      &@      @      &@              @      @      @      �?      @      �?       @              �?      �?      �?      �?                      �?              �?      @      @      @      @      �?      @               @      �?      �?      �?                      �?      @                      �?       @               @              5@      >@      @      8@      @      $@              "@      @      �?       @      �?       @                      �?      @                      ,@      .@      @      &@      @      @      @      @                      @      @              @      @              @      @              @      @              @      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJk�ahG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B@D         
                   @������?�           @�@              S                    �?ް-Z�+�?�           p�@                                    @x�� ���?�            `k@                                "�b@ �O�H�?J            �[@       ������������������������       �        C            �Y@                                03c@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        	       D                   �<@�>���?E             [@       
       #                    �?|�|k6��?:            �U@                                03�@��Sݭg�?            �C@        ������������������������       �                     @               "                  S�-@tk~X��?             B@              !                    �? �o_��?             9@                                 �5@��<b���?             7@                                   �?և���X�?             @                                  �?���Q��?             @                                   .@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                P��+@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   �?      �?             0@        ������������������������       �                     @                                    �?8�Z$���?
             *@                               ���@�8��8��?	             (@        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     &@        $       %                 pf�@�q���?             H@        ������������������������       �                     "@        &       C                 ��1@�99lMt�?            �C@       '       <                    �?     ��?             @@       (       5                    �?�q�q�?             8@       )       4                   �;@�d�����?             3@       *       3                 �[$@�q�q�?
             .@       +       2                   �9@X�Cc�?	             ,@       ,       1                   �6@"pc�
�?             &@        -       .                 �&B@      �?             @        ������������������������       �                     �?        /       0                    0@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        6       ;                    ;@���Q��?             @       7       8                 �̬)@�q�q�?             @        ������������������������       �                     �?        9       :                 @3�/@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        =       B                   �;@      �?              @       >       A                    �?؇���X�?             @       ?       @                 P��%@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        E       F                   �=@����X�?             5@        ������������������������       �                     @        G       J                    �?և���X�?	             ,@        H       I                 ��9$@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        K       R                    C@�z�G��?             $@       L       O                    �?      �?             @        M       N                   �@@      �?             @        ������������������������       �                      @        ������������������������       �                      @        P       Q                 `fV6@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        T       U                    $@8�Uj�?+           0}@        ������������������������       �        
             .@        V       �                    �?��F�?!           @|@        W       x                    �?���Fi�?1            �T@       X       u                   �G@2L�����?'            @Q@       Y       d                     �?f>�cQ�?$            �N@        Z       [                   �:@և���X�?
             ,@        ������������������������       �                     @        \       c                    �?z�G�z�?             $@       ]       b                 p�w@      �?              @       ^       a                 `f�A@؇���X�?             @        _       `                 0C=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        e       h                    0@=QcG��?            �G@        f       g                    '@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        i       j                 ��%@`Ӹ����?            �F@       ������������������������       �                     :@        k       t                    =@�KM�]�?	             3@       l       o                     @؇���X�?             ,@        m       n                 `��,@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        p       s                    �?�C��2(�?             &@        q       r                 `v�0@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        v       w                 ��L@@      �?              @        ������������������������       �                     @        ������������������������       �                     @        y       �                     @և���X�?
             ,@       z       {                   �4@�n_Y�K�?	             *@        ������������������������       �                      @        |       �                 �̾w@���!pc�?             &@       }       ~                    �?z�G�z�?             $@       ������������������������       �                     @               �                 �M@�q�q�?             @        ������������������������       �                      @        �       �                   @K@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ��D:@�V@���?�            w@       �       �                    �?ףp=
�?�            `s@       �       �                 ���!@�ʈD��?�            �r@       �       �                    �?0sS]�?z            �h@        ������������������������       �                     7@        �       �                    �?`���4�?k            �e@       �       �                     @x�g���?i            �e@        ������������������������       �                      @        �       �                 �?�@�{�����?d            �d@       �       �                    �?�:�]��?=            �Y@       �       �                   @@@Hm_!'1�?:            �X@       �       �                   �?@�t����?+             Q@       �       �                 ��@�C��2(�?*            �P@        �       �                    7@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �:@`Jj��?(             O@       �       �                   �5@������?             B@        �       �                   �4@�IєX�?
             1@       ������������������������       �                     $@        �       �                 �1@؇���X�?             @        �       �                  s@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     3@        �       �                 pb@ȵHPS!�?             :@        �       �                 �?$@�q�q�?             "@       �       �                 ��,@؇���X�?             @        ������������������������       �                     @        �       �                   �=@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        
             1@        ������������������������       �                      @        ������������������������       �                     >@        ������������������������       �                     @        �       �                 @3�@�&�5y�?'             O@        �       �                   �D@��.k���?             1@       �       �                   �?@�n_Y�K�?             *@        �       �                    :@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �A@      �?              @       ������������������������       �z�G�z�?             @        ������������������������       ��q�q�?             @        ������������������������       �                     @        �       �                   �0@:	��ʵ�?            �F@        ������������������������       �                     �?        �       �                   �;@fP*L��?             F@        �       �                   �:@�d�����?             3@       �       �                   �3@      �?             0@        �       �                   �2@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     @        �       �                 ��y @HP�s��?             9@       �       �                 ��) @�����H�?             2@       �       �                    ?@�IєX�?             1@       ������������������������       �                     $@        �       �                   �@@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?��9J���?F             Z@       �       �                     @�nkK�?0            @Q@       �       �                     �?��S�ۿ?             �F@        ������������������������       �                     �?        �       �                   �*@t��ճC�?             F@       �       �                   �A@l��\��?             A@       �       �                   �@@H%u��?             9@       �       �                    5@P���Q�?             4@        �       �                   �'@r�q��?             @       �       �                   �1@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     ,@        ������������������������       ����Q��?             @        ������������������������       �                     "@        ������������������������       �                     $@        ������������������������       �                     8@        ������������������������       �                    �A@        �       �                    �?�q�q�?             "@       �       �                 �ܭ2@      �?              @       ������������������������       �                     @        �       �                    :@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    @@����*��?*            �M@        �       �                 `fF<@�d�����?             3@       �       �                   �J@�q�q�?
             (@       �       �                 03k:@�����H�?             "@        ������������������������       �                      @        �       �                   @B@؇���X�?             @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �J@؇���X�?             @       ������������������������       �                     @        �       �                   @>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       	                   D@�G�z�?             D@       �                          �?*;L]n�?             >@       �                           @���>4��?             <@       �       �                  x#J@����X�?             5@        �       �                     �?      �?              @       �       �                   �=@؇���X�?             @       �       �                   �A@z�G�z�?             @        ������������������������       �                      @        �       �                 `f�D@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        �                       ���M@�n_Y�K�?             *@                                  7@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @                              03U@      �?              @       ������������������������       �                     @                                 �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     $@                              ���A@ ��WV�?             :@                                 @ףp=
�?             $@                                 �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             0@        �t�b��     h�h*h-K ��h/��R�(KMKK��h]�B        |@     `p@     �z@     Pp@     �I@      e@      �?     �[@             �Y@      �?      @      �?                      @      I@      M@     �A@      J@      $@      =@      @              @      =@      @      2@      @      2@      @      @       @      @      �?       @               @      �?              �?      �?              �?      �?              �?      �?              �?      �?               @      ,@              @       @      &@      �?      &@      �?                      &@      �?               @                      &@      9@      7@              "@      9@      ,@      2@      ,@      0@       @      ,@      @      $@      @      "@      @      "@       @       @       @              �?       @      �?       @                      �?      @                      @      �?              @               @      @       @      �?      �?              �?      �?              �?      �?                       @       @      @      �?      @      �?      @      �?                      @               @      �?              @              .@      @      @               @      @      �?      @      �?                      @      @      @      @      @       @       @       @                       @      �?      �?              �?      �?              @             `w@     @W@              .@     `w@     �S@     �O@      4@     �K@      ,@      J@      "@       @      @              @       @       @      @       @      @      �?      �?      �?      �?                      �?      @                      �?       @              F@      @      �?      �?      �?                      �?     �E@       @      :@              1@       @      (@       @       @      �?              �?       @              $@      �?      @      �?      @                      �?      @              @              @      @      @                      @       @      @       @      @               @       @      @       @       @      @              @       @       @               @       @       @                       @              �?              �?     ps@      M@     pq@      ?@     q@      <@     �e@      9@      7@             �b@      9@     `b@      9@       @             `a@      9@     �W@       @     �V@       @      N@       @      N@      @       @       @       @                       @      M@      @     �A@      �?      0@      �?      $@              @      �?       @      �?       @                      �?      @              3@              7@      @      @      @      @      �?      @              @      �?       @      �?      �?                       @      1@                       @      >@              @             �F@      1@       @      "@       @      @       @      @       @                      @      @       @      @      �?       @      �?              @     �B@       @              �?     �B@      @      ,@      @      ,@       @      @       @      @                       @      "@                      @      7@       @      0@       @      0@      �?      $@              @      �?              �?      @                      �?      @               @             @Y@      @     �P@      @      E@      @      �?             �D@      @      ?@      @      6@      @      3@      �?      @      �?      @      �?      �?               @      �?       @              ,@              @       @      "@              $@              8@             �A@              @      @      @      @      @              �?      @      �?                      @      �?              @@      ;@      @      ,@      @       @      �?       @               @      �?      @      �?       @              @      @              �?      @              @      �?      �?              �?      �?              ;@      *@      1@      *@      .@      *@      .@      @      @      �?      @      �?      @      �?       @               @      �?              �?       @               @              �?               @      @      �?      @      �?                      @      @      �?      @              @      �?      @                      �?              @       @              $@              9@      �?      "@      �?       @      �?       @                      �?      @              0@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ6ޤhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B@E         �                    �? ��ʀ_�?�           @�@              W                     @�{���2�?X           X�@               <                 `fFJ@|ő����?�            �j@              )                     �? )O7�?]             b@                                  �7@H(���o�?"            �J@        ������������������������       �                      @               
                    �?�q�q�?!            �I@               	                 ���;@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?                                   �?������?            �F@                                `f�A@      �?             (@                               �ܵ<@և���X�?             @        ������������������������       �                     @                                ��>@      �?             @                                 �E@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @               (                 `f�D@���!pc�?            �@@                                 �E@��X��?             <@                                ��$:@���|���?             &@        ������������������������       �                      @                                  `@@�<ݚ�?             "@       ������������������������       �                     @                                  �A@      �?             @        ������������������������       �                      @        ������������������������       �                      @               '                    R@�t����?             1@              &                 `f�;@      �?             0@               !                 ��:@�8��8��?             (@        ������������������������       �                     �?        "       %                    J@�C��2(�?             &@        #       $                   @G@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        *       +                    �?\Ќ=��?;            �V@        ������������������������       �                     >@        ,       /                    �?\#r��?&            �N@        -       .                 hf�2@      �?             @        ������������������������       �                     @        ������������������������       �                     @        0       ;                   �@@�1�`jg�?#            �K@       1       8                   �3@�L���?            �B@       2       7                   �5@г�wY;�?             A@        3       4                   �2@$�q-�?             *@        ������������������������       �                     @        5       6                   �'@      �?              @       ������������������������       �؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     5@        9       :                    8@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     2@        =       L                   �E@��+7��?+            @Q@       >       K                     �?V�a�� �?#             M@       ?       @                    �?PN��T'�?              K@       ������������������������       �                     D@        A       H                    <@և���X�?
             ,@       B       E                    �?      �?              @        C       D                 ���Z@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        F       G                    6@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        I       J                   �B@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        M       R                    �?�eP*L��?             &@       N       O                 @�pX@z�G�z�?             @       ������������������������       �                     @        P       Q                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        S       V                 03oT@r�q��?             @       T       U                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        X       �                    @@��x�?�            `u@       Y       t                    �?R=˄rG�?�            Pu@        Z       s                   @<@     ��?1             T@       [       \                 ��Y@�n_Y�K�?'            @P@        ������������������������       �                     "@        ]       j                    �?h�����?#             L@        ^       g                    �?>���Rp�?             =@       _       `                    �?��s����?             5@        ������������������������       �                      @        a       f                 pF @�	j*D�?             *@       b       c                 ���@"pc�
�?             &@        ������������������������       �                     �?        d       e                 �&B@z�G�z�?             $@       ������������������������       ��<ݚ�?             "@        ������������������������       �                     �?        ������������������������       �                      @        h       i                    �?      �?              @        ������������������������       �                     @        ������������������������       �                     @        k       l                    1@�����H�?             ;@        ������������������������       �                     �?        m       n                    �?$�q-�?             :@        ������������������������       �                     &@        o       r                   @'@�r����?
             .@       p       q                 03�@z�G�z�?             $@        ������������������������       �                     �?        ������������������������       ��<ݚ�?             "@        ������������������������       �                     @        ������������������������       �        
             .@        u       �                    �?T��o��?�            Pp@       v       �                   �;@8�Z$���?�            �n@        w       �                   �:@�W;�E��?G            �Z@       x       �                 �1@�d�$���?C            @Y@        y       �                    �?����e��?            �@@       z       }                   �4@����"�?             =@        {       |                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ~       �                 �?$@�G��l��?             5@              �                    7@�q�q�?             "@       �       �                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �8@      �?             @        ������������������������       �                     �?        �       �                 @33@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�q�q�?             (@       �       �                 ���@؇���X�?             @        ������������������������       �                     @        �       �                   �7@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �6@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ��@      �?             @       ������������������������       �                      @        ������������������������       �                      @        �       �                    �?l��\��?,             Q@       �       �                   �3@�X�<ݺ?$             K@        �       �                   �2@�t����?	             1@       ������������������������       �                     $@        �       �                 �?�@����X�?             @        ������������������������       �                      @        �       �                 `�8"@���Q��?             @       ������������������������       ��q�q�?             @        ������������������������       �                      @        �       �                    �?�?�|�?            �B@        �       �                 pf� @r�q��?             @        �       �                   �8@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     ?@        �       �                   �8@d}h���?             ,@        �       �                   �6@      �?             @       �       �                   �!@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�d�g��?Q            �a@        �       �                    �?���|���?             &@       �       �                    I@�q�q�?             "@       �       �                 `�X!@؇���X�?             @        ������������������������       �                     @        �       �                    A@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                   �B@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?Du9iH��?J             `@       �       �                 �T)D@0{�v��?G            @_@       �       �                   �<@P���Q�?D             ^@        ������������������������       �                    �J@        �       �                 �&B@�qM�R��?(            �P@        ������������������������       �                     4@        �       �                   @@@��E�B��?            �G@        �       �                   �@�E��ӭ�?             2@        ������������������������       �                      @        �       �                   �>@     ��?             0@        �       �                 ���"@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 ��i @      �?              @       �       �                 @3�@�q�q�?             @       �       �                   �?@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �E@XB���?             =@       ������������������������       �        	             1@        �       �                   �F@�8��8��?             (@        �       �                 @3�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        �       �                    >@���Q��?             @       ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     ,@        ������������������������       �                     �?        �       �                     @��>���?b            �c@        �       �                    �?���5��?1            �S@       �       �                    �?�D��?            �H@       ������������������������       �                     9@        �       �                    +@r�q��?             8@        ������������������������       �                     $@        �       �                    �?@4և���?             ,@        �       �                   �@@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     (@        �       �                    @\-��p�?             =@       �       �                 ���`@HP�s��?             9@       �       �                    �?���N8�?             5@       ������������������������       �                     0@        �       �                    �?z�G�z�?             @       �       �                     �?      �?             @        ������������������������       �                      @        �       �                 pV�C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?      �?             @       �       �                    '@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                 @�+@�J�j�?1            �S@        �       �                 pFD @8�Z$���?	             *@        ������������������������       �                      @        ������������������������       �                     &@        �                        �7@"pc�
�?(            �P@        �       �                    $@d��0u��?             >@        �       �                     @      �?              @       ������������������������       �                     @        ������������������������       �                     �?                                  �?"pc�
�?             6@                                 >@�θ�?             *@                                �?�C��2(�?             &@                                  @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @                              8#�1@�����H�?             "@        	      
                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                 �?������?             B@        ������������������������       �                      @                                 @h�����?             <@                              ��T?@�q�q�?             @        ������������������������       �                     �?                                 �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     9@        �t�bh�h*h-K ��h/��R�(KMKK��h]�BP       �|@     �o@     x@     @e@     �Z@     �Z@     @V@     �K@      A@      3@               @      A@      1@      �?      @              @      �?             �@@      (@      "@      @      @      @      @              �?      @      �?      �?              �?      �?                       @      @              8@      "@      3@      "@      @      @       @               @      @              @       @       @       @                       @      .@       @      .@      �?      &@      �?      �?              $@      �?      �?      �?      �?                      �?      "@              @                      �?      @             �K@      B@              >@     �K@      @      @      @              @      @              J@      @      A@      @     �@@      �?      (@      �?      @              @      �?      @      �?      �?              5@              �?       @      �?                       @      2@              2@     �I@      (@      G@       @      G@              D@       @      @      @      @      �?      �?              �?      �?               @      @       @                      @      @      �?      @                      �?      @              @      @      �?      @              @      �?      �?              �?      �?              @      �?       @      �?              �?       @              @             `q@      P@     `q@     �O@     �K@      9@      D@      9@      "@              ?@      9@      @      6@      @      1@               @      @      "@       @      "@              �?       @       @       @      @              �?       @              @      @      @                      @      8@      @              �?      8@       @      &@              *@       @       @       @      �?              @       @      @              .@             �k@      C@      j@      C@     �T@      9@     �T@      3@      4@      *@      2@      &@      @      �?              �?      @              &@      $@      @      @      @      �?              �?      @               @       @              �?       @      �?              �?       @              @      @      �?      @              @      �?      @              @      �?              @      �?              �?      @               @       @       @                       @      O@      @     �I@      @      .@       @      $@              @       @       @              @       @      �?       @       @              B@      �?      @      �?      �?      �?      �?                      �?      @              ?@              &@      @      @      @      @       @               @      @                      �?       @                      @     �_@      *@      @      @      @      @      @      �?      @               @      �?              �?       @                       @      �?      �?              �?      �?              ^@      "@      ]@      "@     �\@      @     �J@             �N@      @      4@             �D@      @      *@      @               @      *@      @      @      �?      @                      �?      @       @      @       @      @      �?              �?      @                      �?       @              <@      �?      1@              &@      �?       @      �?              �?       @              "@               @      @       @      �?               @      @              ,@                      �?     @R@      U@      1@     �N@      *@      B@              9@      *@      &@              $@      *@      �?      �?      �?      �?                      �?      (@              @      9@       @      7@      �?      4@              0@      �?      @      �?      @               @      �?      �?              �?      �?                      �?      �?      @      �?      �?      �?                      �?               @       @       @               @       @              L@      7@       @      &@       @                      &@      K@      (@      3@      &@      �?      @              @      �?              2@      @      $@      @      $@      �?       @      �?       @                      �?       @                       @       @      �?      �?      �?      �?                      �?      @             �A@      �?       @              ;@      �?       @      �?      �?              �?      �?              �?      �?              9@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ��{hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtK�huh*h-K ��h/��R�(KK�h|�B�<         L                    �?^80�B�?�           @�@               =                 �D�H@ �o_��?�            @o@              8                    @�,�:�?_            �d@                                   @P�?�+��?V            �b@        ������������������������       �        !            �J@                                   �?�`���?5            �X@                                  �+@z�G�z�?             D@        ������������������������       �                     @        	                           �?�<ݚ�?             B@        
                           �?�<ݚ�?             2@                                  7@�θ�?             *@        ������������������������       �                     �?                                   �?r�q��?             (@        ������������������������       �                     @                                 S�2@���Q��?             @                                 �<@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?                                   �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @                                   �?�<ݚ�?             2@                                  �?�	j*D�?	             *@                               ���@      �?             (@        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     @               7                   �;@8^s]e�?             M@              2                    �?�\��N��?             C@               !                 ���@`՟�G��?             ?@        ������������������������       �                     @        "       +                    �?��
ц��?             :@       #       $                 P�@������?             1@        ������������������������       �                      @        %       (                 03�!@X�<ݚ�?             "@       &       '                   �8@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        )       *                  �#@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ,       -                    �?�����H�?             "@        ������������������������       �                     @        .       /                    @z�G�z�?             @        ������������������������       �                      @        0       1                    1@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        3       4                    �?؇���X�?             @        ������������������������       �                     @        5       6                 ��6@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     4@        9       <                    @      �?	             0@       :       ;                    =@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        >       K                     @�}#���?0            �T@       ?       @                    �? ���J��?-            �S@        ������������������������       �                     A@        A       B                    �?���7�?             F@       ������������������������       �                     @@        C       J                     �?r�q��?	             (@       D       E                 ���`@      �?              @        ������������������������       �                     @        F       G                    �?      �?             @        ������������������������       �                     �?        H       I                 ���i@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        M       R                    @ӏ�[��?            �|@        N       O                 �Q��?������?             1@        ������������������������       �                     @        P       Q                    @�q�q�?	             (@       ������������������������       �                      @        ������������������������       �                     @        S       �                   @S@&<k����?           �{@       T       �                     �?`���?           �{@        U       �                    @�
I���?;             [@       V       s                    �?$+ޠ�5�?:            @Z@       W       X                   �3@\�CX�?(            �Q@        ������������������������       �                      @        Y       `                    �?2L�����?'            @Q@        Z       _                 p�w@�㙢�c�?             7@       [       \                 ��>@��2(&�?             6@        ������������������������       �                     $@        ]       ^                   �B@      �?             (@        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     �?        a       h                   �B@��<b���?             G@       b       g                   �<@���7�?             6@       c       f                   �>@�X�<ݺ?             2@        d       e                 `f�<@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     @        i       j                 03k:@      �?             8@        ������������������������       �                     @        k       r                   �J@����X�?             5@       l       q                   �G@��
ц��?             *@       m       p                   �F@�z�G��?             $@       n       o                 `f?@և���X�?             @       ������������������������       ����Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        t       u                  x#J@h+�v:�?             A@        ������������������������       �                      @        v       w                 `f�N@     ��?             @@        ������������������������       �                      @        x       }                 Ј�U@r�q��?             8@        y       z                   @G@      �?              @        ������������������������       �                     @        {       |                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ~                        �UcV@     ��?             0@        ������������������������       �                     @        �       �                    �?�eP*L��?             &@        ������������������������       �                     @        �       �                    @؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �T�I@��+�?�            �t@       �       �                 ��y @��XA%��?�            �s@       �       �                    �?p#�����?m            �c@       �       �                     @�"ZN��?d            �b@        ������������������������       �                     @        �       �                 ��) @x�5?,R�?a             b@       �       �                    �?Tri����?`            �a@        �       �                    �?�8��8��?             8@       �       �                   �=@8�Z$���?             *@       �       �                   �<@�<ݚ�?             "@       �       �                 ���@      �?              @        �       �                 ��y@�q�q�?             @        ������������������������       �                     �?        �       �                   �7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             &@        �       �                    1@�S#א��?K            @]@        ������������������������       �                     @        �       �                 @3�@@��xQ�?J            �\@        �       �                   �>@���Q��?             @       �       �                    6@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                   @F@��<nd�?G            @[@       �       �                 �{@�)���Y�?>            �X@        �       �                   �4@$G$n��?            �B@        ������������������������       �                     @        �       �                 �?$@�חF�P�?             ?@       �       �                 ���@�X�<ݺ?             2@        �       �                 ���@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     (@        �       �                   �9@�	j*D�?             *@       �       �                   �5@"pc�
�?             &@       �       �                 �1@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                 �?�@��GEI_�?&            �N@        ������������������������       �                     ?@        �       �                 @3�@�r����?             >@        �       �                   �D@���!pc�?             &@       �       �                    :@z�G�z�?             $@        ������������������������       �                     @        �       �                   �?@����X�?             @        ������������������������       �                     �?        �       �                   �A@r�q��?             @        ������������������������       �                      @        ������������������������       �      �?             @        ������������������������       �                     �?        �       �                    ?@�}�+r��?             3@       ������������������������       �        
             (@        �       �                   �@@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             &@        ������������������������       �                     @        �       �                   �9@�z�G��?	             $@       �       �                    3@      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    !@D���D|�?_            �c@        �       �                    @      �?              @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �9@������?[            �b@        ������������������������       �                    �C@        �       �                    �?��X��?>             \@       �       �                   �:@�Z��L��?&            �Q@        ������������������������       �                      @        �       �                 `f�)@���}<S�?%            @Q@        ������������������������       �                     <@        �       �                    �?�p ��?            �D@        ������������������������       �                      @        �       �                   �*@��-�=��?            �C@        �       �                    =@����X�?	             ,@        ������������������������       �                     �?        �       �                    @@�θ�?             *@        ������������������������       �                     @        �       �                   �F@�z�G��?             $@       �       �                    C@և���X�?             @        ������������������������       �      �?             @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     9@        �       �                    �?��Y��]�?            �D@        ������������������������       �                      @        �       �                   �@@Pa�	�?            �@@       �       �                    ?@��S�ۿ?	             .@       ������������������������       �                     ,@        ������������������������       �                     �?        ������������������������       �                     2@        �       �                    �?X�<ݚ�?             2@       �       �                 ��?P@�q�q�?             (@       �       �                    ;@z�G�z�?             $@        ������������������������       �                     @        �       �                    >@����X�?             @       ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �t�bh�h*h-K ��h/��R�(KK�KK��h]�B0       p{@     q@     �Q@     �f@     �O@      Z@      H@     �Y@             �J@      H@      I@       @      @@              @       @      <@      @      ,@      @      $@      �?               @      $@              @       @      @       @       @       @                       @              �?      �?      @      �?                      @      @      ,@      @      "@      @      "@      @                      "@      �?                      @      D@      2@      4@      2@      ,@      1@              @      ,@      (@      *@      @       @              @      @      �?      @      �?                      @      @      �?      @                      �?      �?       @              @      �?      @               @      �?       @      �?                       @      @      �?      @               @      �?              �?       @              4@              .@      �?      @      �?      @                      �?      "@              @      S@       @      S@              A@       @      E@              @@       @      $@       @      @              @       @       @              �?       @      �?       @                      �?              @      @             w@     @W@      @      *@              @      @       @               @      @             �v@      T@     �v@     �S@     �Q@     �B@      Q@     �B@     �K@      0@               @     �K@      ,@      3@      @      3@      @      $@              "@      @              @      "@                      �?      B@      $@      5@      �?      1@      �?      @      �?      @                      �?      &@              @              .@      "@              @      .@      @      @      @      @      @      @      @       @      @       @              @                      @       @              *@      5@       @              &@      5@               @      &@      *@      @       @      @              @       @               @      @              @      &@              @      @      @      @              �?      @              @      �?              @             `r@     �D@     �q@     �@@      a@      6@      `@      3@      @             @_@      3@     @_@      0@      6@       @      &@       @      @       @      @      �?       @      �?      �?              �?      �?              �?      �?              @                      �?      @              &@             �Y@      ,@              @     �Y@      &@      @       @      �?       @      �?                       @       @              Y@      "@     @V@      "@      @@      @      @              :@      @      1@      �?      @      �?      @                      �?      (@              "@      @      "@       @      @       @               @      @              @                       @     �L@      @      ?@              :@      @       @      @       @       @      @              @       @              �?      @      �?       @              @      �?              �?      2@      �?      (@              @      �?              �?      @              &@                      @      @      @      @      @      @                      @      @             �b@      &@      @       @               @      @             �a@      "@     �C@             �Y@      "@     �O@       @               @     �O@      @      <@             �A@      @               @     �A@      @      $@      @              �?      $@      @      @              @      @      @      @       @       @       @      �?      @              9@              D@      �?       @              @@      �?      ,@      �?      ,@                      �?      2@              $@       @      @       @       @       @              @       @      @       @       @              @       @              @                       @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ?{�hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM+huh*h-K ��h/��R�(KM+��h|�B�J         �                 ��.@�dx<�?�           @�@               5                    �?z����?�            `u@               .                 `ff+@�q�Q�?8             X@              	                     @������?0            �T@                                  �9@ףp=
�?             4@                                   �?���Q��?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                     .@        
                           �?f���M�?%             O@                                  �2@���B���?             :@        ������������������������       �                     @                                   �?�d�����?             3@        ������������������������       �                      @                                `f�@�t����?	             1@                                 �8@      �?             0@        ������������������������       �                     �?                                ���@z�G�z�?             .@        ������������������������       �                     @        ������������������������       �      �?             (@        ������������������������       �                     �?               -                    �?)O���?             B@              ,                    K@     ��?             @@              )                    �?��>4և�?             <@              $                   �;@      �?             8@                                  0@և���X�?             ,@        ������������������������       �                     �?                                pff@�n_Y�K�?
             *@        ������������������������       �                     @               #                  �#@����X�?             @              "                   �!@r�q��?             @                !                    9@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        %       (                    �?ףp=
�?             $@       &       '                   &@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        *       +                   �&@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        /       4                    �?@4և���?             ,@        0       1                 �?�-@؇���X�?             @        ������������������������       �                     @        2       3                   �<@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        6       7                    +@�<p���?�            �n@        ������������������������       �                     @        8       �                    �?��w]j<�?�             n@       9       �                    �?|�9ǣ�?�            �m@       :       ;                     �?@��xQ�?�            �l@        ������������������������       �                     @        <       ]                 �1@�Cc}h��?�             l@        =       Z                    �?��1��?4            �T@       >       Y                   �=@���!���?2            �S@       ?       X                   �<@�S����?%            �L@       @       A                    7@X�;�^o�?$            �K@        ������������������������       �        
             0@        B       C                     @:�&���?            �C@        ������������������������       �                      @        D       E                   �8@��G���?            �B@        ������������������������       �                      @        F       M                    �?؇���X�?            �A@       G       L                    �?�nkK�?             7@       H       I                 ���@�C��2(�?	             &@        ������������������������       �                     @        J       K                   @<@      �?              @       ������������������������       �r�q��?             @        ������������������������       �                      @        ������������������������       �                     (@        N       O                 ��@�q�q�?             (@        ������������������������       �                     �?        P       Q                   �:@���!pc�?             &@        ������������������������       �                      @        R       S                 pf�@�q�q�?             "@        ������������������������       �                      @        T       U                   �;@և���X�?             @        ������������������������       �                     �?        V       W                 �?$@�q�q�?             @       ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     6@        [       \                 ���@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ^       �                    �?,�d�vK�?g            �a@       _       �                 `f�)@���2���?f            �a@       `       g                    �?      �?R             \@        a       f                 �� @؇���X�?             @       b       c                   �<@z�G�z�?             @        ������������������������       �                      @        d       e                    ?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        h       �                   `M@ >�֕�?L            @Z@       i       �                 ���!@X�?٥�?J            �Y@       j       k                 �?�@���;QU�?6            @R@        ������������������������       �                     <@        l       �                   @D@�����H�?!            �F@       m       t                 @3�@�?�'�@�?             C@        n       o                    :@�q�q�?             @        ������������������������       �                     �?        p       q                   �?@���Q��?             @        ������������������������       �                     �?        r       s                   �A@      �?             @        ������������������������       �                      @        ������������������������       �      �?              @        u       ~                 @Q!@     ��?             @@       v       }                 ��i @���}<S�?             7@       w       x                    4@�����?             5@        ������������������������       �                     �?        y       z                    ?@P���Q�?             4@       ������������������������       �                     1@        {       |                   �@@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @               �                   �;@�����H�?             "@       �       �                    6@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     >@        �       �                   �P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 �R,@؇���X�?             <@       �       �                   �;@"pc�
�?             6@        ������������������������       �                     "@        �       �                    �?�	j*D�?             *@        ������������������������       �                     �?        �       �                   �*@      �?
             (@       �       �                    =@�q�q�?             "@        ������������������������       �                     �?        �       �                    @@      �?              @        ������������������������       �                      @        �       �                   �F@�q�q�?             @       �       �                    C@���Q��?             @        ������������������������       �      �?              @        ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �                       ���S@` .�(�?�             w@       �                          @~&���?�            �q@       �       �                    �?�o����?�            �o@        �       �                    �?�t����?'             Q@        ������������������������       �                     D@        �       �                    �?����X�?             <@       �       �                    �?�+e�X�?             9@       �       �                    �?���y4F�?             3@       �       �                    �?r�q��?             2@       �       �                   x5@���!pc�?             &@        �       �                   �2@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    A@      �?              @       �       �                    =@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�q�q�?             @       �       �                   �K@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 pV�C@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �                         R@��;���?w            `g@       �       �                    !@ 9�����?p             f@        ������������������������       �        	             5@        �       �                    �?`%za��?g            `c@        �       �                    �?&ջ�{��?1            @R@       �       �                   �;@�ݜ����?'            �M@        �       �                   �1@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        �       �                   �M@Tt�ó��?"            �H@       �       �                     �?d�
��?             F@       �       �                   �>@     ��?             @@       �       �                 ��$:@@�0�!��?             1@        ������������������������       �                     �?        �       �                    H@      �?
             0@       �       �                   �E@z�G�z�?             $@       �       �                   �?@      �?              @       �       �                 `f�<@      �?             @       ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �        	             .@        �       �                 034@�q�q�?	             (@        ������������������������       �                     @        �       �                   �=@X�<ݚ�?             "@        ������������������������       �                     @        �       �                    >@z�G�z�?             @       �       �                 0�_F@      �?             @        ������������������������       �                      @        ������������������������       �      �?              @        ������������������������       �                     �?        �       �                    R@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    ,@����X�?
             ,@        ������������������������       �                     �?        �       �                    �?�θ�?	             *@       �       �                     @�C��2(�?             &@       ������������������������       �                     "@        �       �                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �8@hP�vCu�?6            �T@        �       �                     @X�<ݚ�?             2@        �       �                    �?؇���X�?             @       �       �                   �4@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    0@���|���?             &@        ������������������������       �                     @        ������������������������       �                     @        �                          �?     ��?+             P@       �                           �?b�2�tk�?             B@       �       �                   �;@���Q��?            �A@        �       �                   �9@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                     @����X�?             <@        ������������������������       �        	             ,@        �       �                    �?և���X�?
             ,@       �       �                    �?      �?              @        �       �                 ��1@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 `fV6@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     <@        ������������������������       �                     &@                                 =@     ��?             @@                                @`Jj��?             ?@                                �?ףp=
�?             4@       ������������������������       �        	             &@                                 �?�<ݚ�?             "@       	      
                ��T?@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?                                 @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     �?              (                   @�1/z��?.            �T@                               �<@�s�c���?,            @S@                                �1@      �?             8@        ������������������������       �                     $@                              `f�n@և���X�?             ,@                                �?�eP*L��?             &@                                �?      �?              @        ������������������������       �                     @                                 �?���Q��?             @        ������������������������       �                     �?                                �5@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @               !                  �G@�&=�w��?            �J@       ������������������������       �                     E@        "      #                   �?"pc�
�?             &@        ������������������������       �                     @        $      '                  �H@���Q��?             @       %      &                ���X@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        )      *                   �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �t�b��     h�h*h-K ��h/��R�(KM+KK��h]�B�       �y@     �r@      p@     �U@     �B@     �M@      8@      M@       @      2@       @      @               @       @      �?              .@      6@      D@      @      5@              @      @      ,@               @      @      (@      @      (@      �?              @      (@              @      @      "@      �?              1@      3@      1@      .@      1@      &@      .@      "@      @       @      �?              @       @              @      @       @      @      �?      �?      �?      �?                      �?      @                      �?      "@      �?       @      �?       @                      �?      �?               @       @       @                       @              @              @      *@      �?      @      �?      @               @      �?       @                      �?      @             `k@      ;@              @     `k@      6@     �j@      6@     �i@      6@      @             @i@      6@     �Q@      &@     �Q@      "@      H@      "@      H@      @      0@              @@      @       @              >@      @               @      >@      @      6@      �?      $@      �?      @              @      �?      @      �?       @              (@               @      @              �?       @      @       @              @      @       @              @      @              �?      @       @      �?       @      @                       @      6@              �?       @      �?                       @     ``@      &@      `@      &@     @Z@      @      @      �?      @      �?       @               @      �?              �?       @               @             �X@      @     �X@      @      Q@      @      <@              D@      @     �@@      @      @       @      �?              @       @              �?      @      �?       @              �?      �?      =@      @      5@       @      3@       @              �?      3@      �?      1@               @      �?              �?       @               @               @      �?      @      �?      @                      �?      @              @              >@              �?      �?              �?      �?              8@      @      2@      @      "@              "@      @              �?      "@      @      @      @              �?      @       @       @              @       @      @       @      �?      �?       @      �?      �?              @              @               @               @              @             `c@     �j@     �a@      b@     @\@     �a@      4@      H@              D@      4@       @      3@      @      .@      @      .@      @       @      @      �?       @      �?                       @      @      �?      @      �?      @                      �?      @              @                      �?      @       @      @       @      @                       @      �?              �?       @               @      �?             @W@     �W@     �T@     �W@              5@     �T@     @R@      @@     �D@      <@      ?@      �?      "@      �?                      "@      ;@      6@      7@      5@      2@      ,@      @      ,@      �?               @      ,@       @       @      �?      @      �?      @      �?      �?               @              @      �?      �?              @      .@              @      @              @      @      @      @              �?      @      �?      @               @      �?      �?              �?      @      �?      @                      �?      @      $@      �?              @      $@      �?      $@              "@      �?      �?              �?      �?               @              I@      @@       @      $@      �?      @      �?      @      �?                      @              �?      @      @              @      @              E@      6@      ,@      6@      ,@      5@      @      �?      @                      �?       @      4@              ,@       @      @       @      @      �?      @              @      �?              �?       @               @      �?              @                      �?      <@              &@              =@      @      =@       @      2@       @      &@              @       @      @      �?      @                      �?      �?      �?              �?      �?              &@                      �?      *@     �Q@       @     @Q@      @      2@              $@      @       @      @      @      @      @              @      @       @      �?               @       @       @                       @      @                      @       @     �I@              E@       @      "@              @       @      @      �?      @              @      �?              �?              @      �?              �?      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ��}whG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B�C         l                     @�K��?�           @�@               	                   �1@$/����?�            Pt@                                    �?ףp=
�?             4@                                   �?�<ݚ�?             "@       ������������������������       �                     @                                ���`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        
             &@        
                           �?��*��?�            s@                                  �;@T��,��?E            @Y@                                   �?l��\��?             A@                               ��*@P���Q�?             4@                                  �'@؇���X�?             @        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     *@                                  �8@؇���X�?             ,@       ������������������������       �                     (@        ������������������������       �                      @        ������������������������       �        2            �P@                                   :@��[�8��?p            �i@                                   4@���7�?             6@                                  �2@      �?              @        ������������������������       �                     @                                    �?      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     ,@               7                 `fF:@LfK!��?c            �f@               6                    �?p`q�q��?+            �S@               %                    �?�:�^���?*            �S@        !       $                    �?և���X�?             @       "       #                 ���,@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        &       5                   �M@����Q8�?'            �Q@       '       (                 `f�)@hA� �?&            �Q@        ������������������������       �                     <@        )       .                   �<@@4և���?             E@        *       -                   �*@�q�q�?             @        +       ,                   �;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        /       4                   �*@������?             B@        0       1                   @D@$�q-�?             *@        ������������������������       �                     @        2       3                   �F@؇���X�?             @        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     7@        ������������������������       �                     �?        ������������������������       �                     �?        8       ;                   �;@�ԇ���?8            �Y@        9       :                    �?���|���?             &@       ������������������������       �                     @        ������������������������       �                     @        <       E                   �>@�)
;&��?4             W@        =       D                   �<@r�q��?             8@       >       ?                    �?���y4F�?             3@        ������������������������       �                     @        @       C                   �>@������?             .@        A       B                 `fF<@և���X�?             @        ������������������������       ����Q��?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        F       S                    �?�v:���?%             Q@        G       J                   �A@�q�����?             9@        H       I                    �?���!pc�?             &@        ������������������������       �                      @        ������������������������       �                     @        K       R                    �?X�Cc�?             ,@       L       O                    �?�eP*L��?             &@        M       N                   �B@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        P       Q                   �H@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        T       a                    @@^����?            �E@        U       \                   �J@      �?
             2@       V       [                    �?���!pc�?             &@       W       X                 `f�;@z�G�z�?             $@       ������������������������       �                     @        Y       Z                   �=@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ]       ^                 `fF<@؇���X�?             @        ������������������������       �                     @        _       `                   @>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        b       c                 ��9L@H%u��?             9@        ������������������������       �                     $@        d       i                    �?z�G�z�?	             .@       e       h                    �?8�Z$���?             *@       f       g                 03�M@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        j       k                 ���Y@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        m                        ��Y7@����G��?�            0x@       n       �                    �?f���]�?�            �s@        o       �                 ��.@N֩	%��?4            @V@       p       q                 P�*@.}Z*�?)            �Q@        ������������������������       �                     @        r       �                    �?     8�?%             P@       s       |                    �?TV����?#            �M@        t       {                    �?l��
I��?             ;@       u       z                 pF @�㙢�c�?             7@       v       y                 ���@�����?             5@        w       x                 0��@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �                      @        ������������������������       �                     @        }       �                   �7@     ��?             @@        ~       �                   �5@      �?             @              �                 ���@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   @<@؇���X�?             <@       �       �                   �:@���y4F�?             3@        ������������������������       �                     @        �       �                    �?������?
             .@        �       �                 ���@      �?             @        ������������������������       �                     �?        ������������������������       ����Q��?             @        ������������������������       ������H�?             "@        ������������������������       �                     "@        �       �                    +@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ��6@r�q��?             2@       �       �                    �?�θ�?             *@        �       �                   x4@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?z�G�z�?             $@       �       �                    �?�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?��m��?�            �l@        �       �                   �K@Rg��J��?#            �H@       �       �                    �?z�J��?"            �G@       �       �                    @����e��?            �@@       �       �                   @D@      �?             @@       �       �                    �?���Q��?             >@       �       �                   �@@�f7�z�?             =@       �       �                    3@��>4և�?             <@        �       �                    0@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �4@��H�}�?             9@        ������������������������       �                     @        �       �                 ��1@8�A�0��?             6@       �       �                 �̬)@      �?             2@       �       �                   �>@�n_Y�K�?             *@       �       �                 @3�@���!pc�?
             &@       �       �                    �?      �?             @       �       �                 ���@���Q��?             @        ������������������������       �                     �?        �       �                 �&B@      �?             @        ������������������������       �                     �?        �       �                   �8@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    9@z�G�z�?             @        ������������������������       �                      @        �       �                    ;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                 ���4@d}h���?
             ,@       �       �                 P��%@�C��2(�?             &@        �       �                    �?z�G�z�?             @        ������������������������       �                      @        �       �                    @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 @3�@d��ϸ�?v            `f@       �       �                 �?�@�?a/��?>            �T@       �       �                 �{@�7�QJW�?8            �R@       �       �                    A@����|e�?&             K@       �       �                    7@�q�q�?            �C@        �       �                 �?$@�X�<ݺ?             2@       ������������������������       �                     (@        �       �                 �1@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?և���X�?             5@       �       �                   �;@�\��N��?             3@       �       �                    :@�n_Y�K�?             *@       �       �                 @33@X�<ݚ�?             "@        ������������������������       �                     @        �       �                   �8@r�q��?             @        �       �                   �@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    >@�q�q�?             @       �       �                 pf�@z�G�z�?             @       ������������������������       �                     @        �       �                 �?$@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     .@        ������������������������       �                     5@        �       �                    :@      �?              @        ������������������������       �                     �?        �       �                   �?@����X�?             @        ������������������������       �                     �?        �       �                   �A@�q�q�?             @        ������������������������       ��q�q�?             @        ������������������������       ��q�q�?             @        �       �                    &@      �?8             X@        �       �                    @      �?              @        ������������������������       �                     @        ������������������������       �                     @        �       �                    ;@�|���?4             V@        ������������������������       �                    �@@        �       �                    �? �Jj�G�?            �K@       �       �                   �<@��Y��]�?            �D@        �       �                 ��) @��S�ۿ?
             .@       ������������������������       �                     $@        �       �                 �̜!@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     :@        ������������������������       �                     ,@                                 �?(N:!���?&            �Q@                                 >@��S���?             .@                             �T)D@z�G�z�?             $@        ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                     @                                 �? �Jj�G�?            �K@        ������������������������       �        
             1@        	                      ��p@@P�Lt�<�?             C@        
                         @�8��8��?	             (@                                 @�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     :@        �t�bh�h*h-K ��h/��R�(KMKK��h]�B�       @|@     @p@     �d@      d@       @      2@       @      @              @       @      �?              �?       @                      &@     `d@     �a@      @     �X@      @      ?@      �?      3@      �?      @              @      �?      �?              *@       @      (@              (@       @                     �P@      d@      F@      5@      �?      @      �?      @              @      �?      �?               @      �?      ,@             `a@     �E@      R@      @     �Q@      @      @      @      �?      @              @      �?              @             �P@      @     �P@      @      <@             �C@      @      @       @      �?       @      �?                       @      @             �A@      �?      (@      �?      @              @      �?      @      �?      @              7@                      �?      �?             �P@      B@      @      @              @      @             �O@      =@      4@      @      .@      @      @              &@      @      @      @      @       @               @       @              @             �E@      9@      (@      *@      @       @               @      @              "@      @      @      @      @       @               @      @              �?      @              @      �?              @              ?@      (@      "@      "@      @       @       @       @              @       @       @       @                       @      �?              @      �?      @              �?      �?              �?      �?              6@      @      $@              (@      @      &@       @      @       @               @      @              @              �?      �?      �?                      �?     �q@      Y@      l@      W@     �G@      E@      F@      ;@      @             �B@      ;@     �@@      :@       @      3@      @      3@       @      3@       @       @               @       @                      &@       @              @              9@      @      �?      @      �?      �?              �?      �?                       @      8@      @      .@      @      @              &@      @      @      @      �?               @      @       @      �?      "@              @      �?              �?      @              @      .@      @      $@      �?       @               @      �?               @       @      �?       @      �?                       @      �?                      @     @f@      I@      7@      :@      7@      8@      4@      *@      4@      (@      2@      (@      1@      (@      1@      &@      �?       @      �?                       @      0@      "@      @              *@      "@      "@      "@       @      @       @      @      @      @       @      @              �?       @       @      �?              �?       @      �?                       @      �?              @                       @      �?      @               @      �?       @      �?                       @      @                      �?      �?               @                      �?      @      &@      �?      $@      �?      @               @      �?       @      �?                       @              @       @      �?       @                      �?               @     `c@      8@     @P@      2@      O@      *@     �D@      *@      :@      *@      1@      �?      (@              @      �?              �?      @              "@      (@      "@      $@      @       @      @      @              @      @      �?      �?      �?              �?      �?              @                      @      @       @      @      �?      @              �?      �?              �?      �?                      �?               @      .@              5@              @      @      �?               @      @              �?       @      @      �?       @      �?       @     �V@      @      @      @      @                      @     �U@      �?     �@@              K@      �?      D@      �?      ,@      �?      $@              @      �?              �?      @              :@              ,@              O@       @       @      @       @       @      @              @       @              @      K@      �?      1@             �B@      �?      &@      �?       @      �?       @                      �?      "@              :@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�,�hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMOhuh*h-K ��h/��R�(KMO��h|�B�S         p                    �?\H�l�?�           @�@                                   �?�-��T��?�            �o@                                  �4@�y��*�?#             M@                                033.@      �?             4@                                  �"@      �?              @        ������������������������       �                     �?                                  �-@����X�?             @        ������������������������       �                      @        	       
                    0@���Q��?             @        ������������������������       �                     �?                                  �1@      �?             @                                Su*@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     (@                                    @�}�+r��?             C@       ������������������������       �                     <@                                   @z�G�z�?             $@                                  �?      �?              @                                H�%@      �?             @        ������������������������       �                     @        ������������������������       �                     �?                                 S�2@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @               o                    @`�'�?w            �h@              T                    �?�z�G��?s            �g@              /                    �?���!pc�?H            @^@               .                    �?r�q��?             >@               !                 ���@���B���?             :@        ������������������������       �                     �?        "       #                   �2@�J�4�?             9@        ������������������������       �                     @        $       %                     @��s����?             5@        ������������������������       �                     @        &       -                 pF @������?             1@       '       (                   �5@�r����?
             .@        ������������������������       �                     �?        )       *                    9@@4և���?	             ,@        ������������������������       �                     �?        +       ,                 �&B@$�q-�?             *@       ������������������������       �ףp=
�?             $@        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        0       S                     @�	j*D�?6            �V@       1       H                    �?l�Ӑ���?4            �U@       2       7                     @L
�q��?%            �M@       3       6                   �9@     ��?             @@        4       5                     �?      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     :@        8       9                 pf�@��}*_��?             ;@        ������������������������       �                     @        :       =                   �9@��+7��?             7@        ;       <                    4@$�q-�?             *@        ������������������������       �                     �?        ������������������������       �                     (@        >       A                 �?�@      �?             $@        ?       @                   �@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        B       C                   �;@�q�q�?             @        ������������������������       �                     @        D       E                    =@�q�q�?             @        ������������������������       �                     �?        F       G                   &@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        I       J                 ���.@����X�?             <@        ������������������������       �                     @        K       N                   �;@r�q��?             8@        L       M                    9@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        O       P                     @�}�+r��?	             3@       ������������������������       �                     (@        Q       R                 03�1@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        U       Z                     @�LQ�1	�?+            @Q@       V       W                 ���`@�FVQ&�?            �@@       ������������������������       �                     :@        X       Y                 Ъ�c@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        [       h                   �;@b�2�tk�?             B@       \       _                    �?և���X�?             5@        ]       ^                 P��%@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        `       a                    �?     ��?
             0@        ������������������������       �                     @        b       c                    @�z�G��?             $@        ������������������������       �                     @        d       g                 ��T?@      �?             @       e       f                    ,@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        i       n                    �?�r����?             .@       j       m                     @z�G�z�?             $@       k       l                 03S1@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        q       �                     �?
"����?$           �|@        r       s                    &@��+7��?;             W@        ������������������������       �                     @        t       �                    �?��~l�?9            @V@       u       ~                    �?`��:�?(            �N@        v       w                    ?@8�Z$���?
             *@        ������������������������       �                      @        x       }                 ڪ�q@���Q��?             @       y       |                    �?      �?             @       z       {                    A@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?               �                   �>@�q�q�?             H@       �       �                   @>@���!pc�?            �@@       �       �                   �Q@z�G�z�?             >@       �       �                   �F@؇���X�?             <@       �       �                 ��I/@      �?
             0@        ������������������������       �                     @        �       �                    @@���Q��?             $@        ������������������������       �                     @        �       �                 03k:@և���X�?             @        ������������������������       �                     @        ������������������������       �      �?             @        ������������������������       �                     (@        ������������������������       �                      @        ������������������������       �                     @        �       �                 `f�D@��S�ۿ?             .@       �       �                   �A@؇���X�?             @       ������������������������       �                     @        �       �                   @B@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ���X@��X��?             <@       �       �                  x#J@�û��|�?             7@        ������������������������       �                     @        �       �                   �D@�\��N��?             3@       �       �                 `f�N@�n_Y�K�?             *@        ������������������������       �                     @        �       �                 0w�U@      �?              @       ������������������������       �                     @        ������������������������       �                     @        �       �                 �UwR@r�q��?             @        ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �                           $@�}�J;��?�            �v@       �       �                   @@�P�I[��?�            �i@        �       �                    �?8�Z$���?:            �V@        �       �                    �?�<ݚ�?             ;@       �       �                   �7@�+e�X�?             9@        �       �                    5@X�<ݚ�?             "@        �       �                 �{@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                 ���@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    =@      �?             0@       �       �                   �:@�C��2(�?             &@        ������������������������       �                     �?        �       �                 ���@ףp=
�?             $@        ������������������������       �                     @        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?      �?*             P@        ������������������������       �        
             .@        �       �                     @ZՏ�m|�?             �H@        ������������������������       �                     @        �       �                   �=@"pc�
�?             F@       �       �                 �?$@�	j*D�?             :@       �       �                    �?�<ݚ�?             2@       �       �                    7@z�G�z�?             .@        ������������������������       �                      @        �       �                   �8@և���X�?             @        ������������������������       �                     �?        �       �                 @33@�q�q�?             @        ������������������������       �                     �?        �       �                 pf�@z�G�z�?             @        ������������������������       �                      @        �       �                    ;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        �       �                 ��@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �6@      �?              @        ������������������������       �                      @        �       �                   �9@�q�q�?             @        ������������������������       �                      @        �       �                   �;@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        	             2@        �       �                ��k @l�b�G��?J            �\@        ������������������������       �                     �?        �       �                    �? (��?I            @\@       �       �                   �3@��Wv��?E             [@        �       �                   �0@؇���X�?
             ,@        �       �                 pFD!@z�G�z�?             @       ������������������������       ��q�q�?             @        ������������������������       �                      @        �       �                    2@�����H�?             "@        ������������������������       �                     @        �       �                 �?�@z�G�z�?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        �       �                 �?�@��ɹ?;            �W@        �       �                 ��@��?^�k�?            �A@        ������������������������       �                     @        �       �                   �<@XB���?             =@       ������������������������       �                     1@        �       �                    �?�8��8��?             (@        �       �                    ?@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 @3�@ ,��-�?$            �M@        �       �                   �A@r�q��?             @        ������������������������       �                     @        ������������������������       �      �?              @        �       �                   @:@ �h�7W�?             �J@        ������������������������       �                     1@        �       �                 ��) @�8��8��?             B@       �       �                    ?@P���Q�?             4@       ������������������������       �                     *@        �       �                   �@@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �>@      �?	             0@       �       �                   �<@z�G�z�?             $@       �       �                 �̜!@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ���"@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @              6                ��Y7@     ��?e             d@             )                   �?R�L=��?:            @X@                                !@��2(&�?'            �P@        ������������������������       �                     �?              "                    @�?�<��?&            @P@                               �;@���c���?             J@                                 &@P���Q�?             4@                                �5@r�q��?             @        	      
                  �1@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     ,@                              ��\+@     ��?             @@                               �A@\-��p�?             =@                             `fF)@     ��?	             0@        ������������������������       �                     @                                �*@���!pc�?             &@                                =@�q�q�?             "@        ������������������������       �                     �?                                 @@      �?              @        ������������������������       �                     @        ������������������������       �      �?             @        ������������������������       �                      @                                 �?$�q-�?             *@        ������������������������       �                      @                                 L@�C��2(�?             &@       ������������������������       �                     @                                �P@      �?             @        ������������������������       �                     �?        ������������������������       �                     @               !                  �B@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        #      (                   �?$�q-�?             *@       $      '                   �?      �?              @        %      &                  �2@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        *      +                ��&@f���M�?             ?@        ������������������������       �                     @        ,      5                   @����X�?             <@       -      .                   �?l��
I��?             ;@        ������������������������       �                     �?        /      0                   #@R�}e�.�?             :@        ������������������������       �                     @        1      2                   �?�����?             5@       ������������������������       �                     1@        3      4                   �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        7      8                ��T?@�[|x��?+            �O@       ������������������������       �                    �A@        9      >                   �?�>4և��?             <@        :      =                pV�C@z�G�z�?             @       ;      <                   �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ?      H                   �?�㙢�c�?             7@        @      A                   *@և���X�?             @        ������������������������       �                     �?        B      C                    @�q�q�?             @        ������������������������       �                      @        D      E                   ;@      �?             @        ������������������������       �                     �?        F      G                   >@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        I      J                   �?      �?             0@        ������������������������       �                     @        K      N                   @ףp=
�?             $@        L      M                   @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �t�bh�h*h-K ��h/��R�(KMOKK��h]�B�       �|@     �o@     �Q@      g@      @     �I@      @      .@      @      @              �?      @       @       @              @       @              �?      @      �?       @      �?              �?       @              �?                      (@       @      B@              <@       @       @       @      @      �?      @              @      �?              �?      @      �?                      @               @      P@     �`@     �L@     �`@     �@@      V@      @      9@      @      5@      �?              @      5@              @      @      1@              @      @      *@       @      *@      �?              �?      *@              �?      �?      (@      �?      "@              @       @                      @      <@     �O@      <@     �M@      4@     �C@      @      =@      @      @              @      @                      :@      1@      $@              @      1@      @      (@      �?              �?      (@              @      @      @      �?              �?      @               @      @              @       @      �?      �?              �?      �?      �?                      �?       @      4@      @              @      4@      @       @               @      @              �?      2@              (@      �?      @              @      �?                      @      8@     �F@       @      ?@              :@       @      @       @                      @      6@      ,@      "@      (@       @      @       @                      @      @      "@              @      @      @      @              @      @      @      �?      @                      �?               @      *@       @       @       @      @       @      @                       @      @              @              @              x@     �Q@      Q@      8@              @      Q@      5@     �H@      (@      &@       @       @              @       @      @      �?       @      �?              �?       @              �?                      �?      C@      $@      8@      "@      8@      @      8@      @      (@      @      @              @      @      @              @      @              @      @      �?      (@                       @              @      ,@      �?      @      �?      @              �?      �?              �?      �?               @              3@      "@      ,@      "@      @              $@      "@      @       @              @      @      @      @                      @      @      �?      @               @      �?              �?       @              @             �s@     �G@     �f@      6@     @S@      ,@      5@      @      3@      @      @      @       @      @       @                      @       @       @               @       @              .@      �?      $@      �?      �?              "@      �?      @              @      �?      @               @              L@       @      .@             �D@       @      @              B@       @      2@       @      ,@      @      (@      @       @              @      @              �?      @       @              �?      @      �?       @               @      �?      �?              �?      �?       @      �?       @                      �?      @      @               @      @       @       @               @       @               @       @              2@             �Z@       @              �?     �Z@      @     @Y@      @      (@       @      @      �?       @      �?       @               @      �?      @              @      �?       @               @      �?     @V@      @      A@      �?      @              <@      �?      1@              &@      �?      @      �?              �?      @              @             �K@      @      @      �?      @              �?      �?      I@      @      1@             �@@      @      3@      �?      *@              @      �?              �?      @              ,@       @       @       @      @      �?              �?      @               @      �?       @                      �?      @              @             �`@      9@     @S@      4@     �L@      "@              �?     �L@       @     �F@      @      3@      �?      @      �?       @      �?       @                      �?      @              ,@              :@      @      9@      @      *@      @      @               @      @      @      @              �?      @       @      @               @       @       @              (@      �?       @              $@      �?      @              @      �?              �?      @              �?       @               @      �?              (@      �?      @      �?       @      �?       @                      �?      @              @              4@      &@              @      4@       @      3@       @              �?      3@      @              @      3@       @      1@               @       @               @       @              �?              M@      @     �A@              7@      @      @      �?       @      �?       @                      �?       @              3@      @      @      @              �?      @       @       @               @       @              �?       @      �?       @                      �?      .@      �?      @              "@      �?       @      �?              �?       @              @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�%\hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B@F                            @^80�B�?�           @�@              �                  x#J@�5j��?�           8�@              J                    �?�q�q�?f           �@               )                 `f�$@R�W�I��?x            �h@                                   �?��o	��?$             M@                                   9@�E��ӭ�?             2@        ������������������������       �                     @                                `f�@X�Cc�?	             ,@       	       
                    �?      �?             (@        ������������������������       �                     �?                                 ��@���!pc�?             &@        ������������������������       �                     �?                                ���@z�G�z�?             $@        ������������������������       �                     �?        ������������������������       ��<ݚ�?             "@        ������������������������       �                      @                                ���@��Q��?             D@        ������������������������       �                     @               $                   �;@�E��ӭ�?             B@              #                  �M$@      �?             8@              "                   �9@և���X�?             5@              !                   �6@�t����?
             1@                                   �?      �?             $@                                  5@X�<ݚ�?             "@                                  3@      �?              @                                  0@      �?             @        ������������������������       �                     �?                                ��!@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        %       &                 `�X!@�8��8��?             (@       ������������������������       �                     @        '       (                 `�("@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        *       +                     @��+7��?T            @a@       ������������������������       �        /             S@        ,       I                 ��Y7@�P�*�?%             O@       -       H                 `v�5@�ՙ/�?             E@       .       7                    �?D�n�3�?             C@        /       0                 �?�-@X�<ݚ�?             "@        ������������������������       �                     @        1       6                    �?z�G�z�?             @       2       3                    -@      �?             @        ������������������������       �                      @        4       5                   �<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        8       E                    �?����"�?             =@       9       :                    �?      �?
             0@        ������������������������       �                     @        ;       <                    �?�q�q�?             (@        ������������������������       �                     �?        =       D                   �=@���|���?             &@       >       C                    ;@և���X�?             @       ?       B                    �?      �?             @       @       A                    9@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        F       G                 ���4@�θ�?             *@       ������������������������       �                     $@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        
             4@        K       j                     �?�&�ѩ��?�            �w@        L       M                   �;@�	j*D�?#             J@        ������������������������       �                     �?        N       S                    �?�t����?"            �I@        O       P                    ?@�<ݚ�?             "@       ������������������������       �                     @        Q       R                    A@      �?             @        ������������������������       �                      @        ������������������������       �                      @        T       c                   �>@��i#[�?             E@       U       V                   �9@      �?             8@        ������������������������       �                     @        W       X                   �<@�q�q�?             2@        ������������������������       �                     @        Y       Z                    @@      �?
             (@        ������������������������       �                      @        [       \                 03k:@���Q��?	             $@        ������������������������       �                      @        ]       b                 `fF<@      �?              @       ^       a                   �K@և���X�?             @        _       `                   @G@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        d       i                   �=@�X�<ݺ?             2@        e       f                   �A@؇���X�?             @        ������������������������       �                     @        g       h                 ��yC@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        k       �                 �?�@�&��?�            Pt@        l       {                    �?�=|+g��?H            @\@        m       n                 03S@��+7��?             7@        ������������������������       �                      @        o       p                   �7@����X�?             5@        ������������������������       �                      @        q       r                 ���@���y4F�?             3@        ������������������������       �                     @        s       v                   @@�q�q�?
             (@       t       u                   @<@      �?              @       ������������������������       �      �?             @        ������������������������       �                      @        w       x                   �<@      �?             @        ������������������������       �                      @        y       z                    ?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        |       �                    �?`Ӹ����?8            �V@       }       ~                   �:@��+��<�?5            �U@        ������������������������       �                    �B@               �                 ��@��<D�m�?"            �H@        ������������������������       �                     8@        �       �                    �?H%u��?             9@        ������������������������       �                     �?        �       �                   �;@      �?             8@        ������������������������       �                     �?        �       �                   �@���}<S�?             7@        �       �                 �&B@�<ݚ�?             "@       �       �                   �>@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    D@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        
             ,@        �       �                 ��@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�iʫ{�?�            �j@        �       �                     @�����?             3@        �       �                    �?      �?              @       �       �                   �<@؇���X�?             @        �       �                 ���,@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                 =
�@���|���?             &@        ������������������������       �                      @        �       �                    '@�<ݚ�?             "@        ������������������������       �                      @        �       �                    3@����X�?             @        ������������������������       �                     �?        �       �                    �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    )@��|���?x             h@        �       �                     @�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        �       �                 @3�@�1j�P�?p            �f@        �       �                    �?�eP*L��?             &@       �       �                   �4@�q�q�?             "@        ������������������������       �                      @        �       �                    :@և���X�?             @        ������������������������       �                      @        �       �                   �?@z�G�z�?             @        ������������������������       �                      @        �       �                    C@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?`ۘV�?i            @e@        �       �                   `3@      �?              @       ������������������������       �                     @        �       �                 03�7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�>����?c            @d@       �       �                   �*@�C��2(�?M            @^@       �       �                 ��) @�+�$f��?A            �X@        �       �                   �3@�X�<ݺ?             B@        �       �                   �1@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        �       �                    ?@Pa�	�?            �@@       ������������������������       �                     5@        �       �                   �@@�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        �       �                    �?���-T��?)             O@       �       �                     @f>�cQ�?(            �N@       �       �                 `fF)@��-�=��?            �C@        ������������������������       �        	             1@        �       �                   �:@"pc�
�?             6@       ������������������������       �                     *@        �       �                   @B@X�<ݚ�?             "@        �       �                    =@z�G�z�?             @        ������������������������       �                      @        �       �                    @@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   �8@�GN�z�?             6@        ������������������������       �                      @        �       �                   �>@X�Cc�?
             ,@       �       �                   �;@      �?              @        ������������������������       �                      @        �       �                   �<@      �?             @       �       �                 �̜!@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                 ���"@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     7@        �       �                     @��Y��]�?            �D@        �       �                    :@�}�+r��?	             3@       �       �                   �7@�C��2(�?             &@        ������������������������       �                      @        �       �                   �<@�����H�?             "@        ������������������������       �                     @        �       �                   �@@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     6@        �                           �?���΍L�?@            �Z@       �       �                 `��M@*S%��?;            �X@        ������������������������       �                     7@        �                         �B@|�i���?0             S@       �       �                    �? s�n_Y�?             J@       �       �                   �A@��hJ,�?             A@       �       �                    �? 	��p�?             =@       ������������������������       �                     6@        �       �                 p�w@����X�?             @       �       �                 ��V\@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                 0w�Z@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �                          <@�q�q�?
             2@       �       �                    3@���Q��?             $@        ������������������������       �                     @        �                        0U�o@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @                              ��Q@      �?             8@        ������������������������       �                     @                                 �?և���X�?             5@       ������������������������       �        	             &@              
                @�pX@ףp=
�?             $@             	                Ј�U@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @                                 >@և���X�?             @                             ��?P@z�G�z�?             @                                ;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @                                 @�C��2(�?            �@@                                �?z�G�z�?             .@        ������������������������       �                      @                              ��T?@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     2@        �t�b� (     h�h*h-K ��h/��R�(KMKK��h]�B�       p{@     q@     �y@     �p@     �w@     �g@     �P@      `@      ?@      ;@      @      *@              @      @      "@      @      "@              �?      @       @      �?               @       @              �?       @      @       @              :@      ,@              @      :@      $@      .@      "@      (@      "@      (@      @      @      @      @      @      @      @      @      @      �?               @      @       @                      @       @                      �?              �?      @                      @      @              &@      �?      @              @      �?              �?      @              B@     �Y@              S@      B@      :@      0@      :@      0@      6@      @      @      @              �?      @      �?      @               @      �?      �?      �?                      �?              �?      &@      2@       @       @              @       @      @      �?              @      @      @      @      @      �?       @      �?              �?       @              �?                      @      @              @      $@              $@      @                      @      4@             �s@      O@      B@      0@              �?      B@      .@      @       @      @               @       @               @       @              =@      *@      (@      (@      @              @      (@              @      @      @       @              @      @               @      @      @      @      @      �?      @      �?                      @      @                      �?      1@      �?      @      �?      @              @      �?              �?      @              &@             pq@      G@     �Y@      $@      1@      @       @              .@      @               @      .@      @      @               @      @      @      @      @      @       @              @      �?       @              �?      �?              �?      �?             �U@      @     �T@      @     �B@              G@      @      8@              6@      @      �?              5@      @              �?      5@       @      @       @      @      �?              �?      @               @      �?              �?       @              ,@              @      �?      @                      �?      f@      B@      *@      @      @       @      @      �?      �?      �?              �?      �?              @                      �?      @      @               @      @       @       @              @       @              �?      @      �?              �?      @             `d@      >@      �?      &@              &@      �?             @d@      3@      @      @      @      @               @      @      @       @              �?      @               @      �?       @      �?                       @       @             �c@      *@      @      �?      @              �?      �?              �?      �?             �b@      (@     �[@      &@     �U@      &@      A@       @       @      �?      �?              �?      �?      @@      �?      5@              &@      �?              �?      &@             �J@      "@      J@      "@     �A@      @      1@              2@      @      *@              @      @      �?      @               @      �?       @      �?                       @      @              1@      @       @              "@      @      @      @               @      @      @       @       @               @       @              �?      �?      �?                      �?      @              �?              7@              D@      �?      2@      �?      $@      �?       @               @      �?      @              @      �?              �?      @               @              6@              ;@     �S@      7@      S@              7@      7@     �J@      &@     �D@      @      =@       @      ;@              6@       @      @       @       @               @       @                      @      @       @      @                       @      @      (@      @      @              @      @      �?      @                      �?               @      (@      (@      @              "@      (@              &@      "@      �?      @      �?      @                      �?      @              @      @      @      �?       @      �?              �?       @               @                       @      >@      @      (@      @       @              @      @      @                      @      2@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ2�hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMChuh*h-K ��h/��R�(KMC��h|�B�P         v                  �#@�Qc�!�?�           @�@               -                    �?6�����?�            �q@                                   �?�m����?'            �M@                                �Y�@�q�q�?             8@        ������������������������       �                      @                                Ь* @���!pc�?             6@              
                   �5@���N8�?             5@               	                   �2@      �?             @       ������������������������       �                     @        ������������������������       �                     @                                   9@�r����?
             .@        ������������������������       �                      @                                0��@8�Z$���?	             *@        ������������������������       �                     @                                 ��@z�G�z�?             $@        ������������������������       �                     �?                                ���@�����H�?             "@        ������������������������       �                     �?                                �&B@      �?              @       ������������������������       �؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     �?                                ���@���Q��?            �A@        ������������������������       �                     @               ,                    �?�c�Α�?             =@              +                    �?���B���?             :@              *                    K@�E��ӭ�?             2@                                  5@������?             1@        ������������������������       �                     @               )                 `��!@�	j*D�?             *@              (                 `�X!@���Q��?             $@               '                 @3�@      �?              @       !       "                 ��@���Q��?             @        ������������������������       �                      @        #       $                   �6@�q�q�?             @        ������������������������       �                     �?        %       &                   �8@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        .       e                 @� @���Lͩ�?�             l@       /       d                   @@@<2r�Y�?z             h@       0       Y                 �{@tX�}}��?^            �b@       1       V                   �?@��� ��?9            @W@       2       3                    7@�����H�?7            �V@        ������������������������       �                     <@        4       5                     @�חF�P�?'             O@        ������������������������       �                     $@        6       =                 ��@���B���?!             J@        7       8                   �8@���Q��?             @        ������������������������       �                      @        9       :                 P��@�q�q�?             @        ������������������������       �                     �?        ;       <                    :@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        >       S                    �?��0{9�?            �G@       ?       @                   �:@X�EQ]N�?            �E@        ������������������������       �                     "@        A       P                 �?$@��hJ,�?             A@       B       I                  s�@      �?             @@        C       H                    =@      �?             0@       D       G                 �Y�@@4և���?	             ,@       E       F                 ���@      �?              @        ������������������������       �                     �?        ������������������������       �؇���X�?             @        ������������������������       �                     @        ������������������������       �                      @        J       O                    >@     ��?             0@       K       N                 ��@�θ�?	             *@       L       M                   �<@z�G�z�?             $@       ������������������������       ������H�?             "@        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     @        Q       R                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        T       U                 �&B@      �?             @        ������������������������       �                      @        ������������������������       �                      @        W       X                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        Z       [                    �?�8���?%             M@        ������������������������       �                     �?        \       ]                    1@���U�?$            �L@        ������������������������       �                     �?        ^       _                 @3�@�h����?#             L@        ������������������������       �                     7@        `       c                 ��Y @Pa�	�?            �@@       a       b                    ?@      �?             @@       ������������������������       �                     ?@        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     E@        f       u                    �?     ��?             @@       g       h                   �9@�r����?             >@        ������������������������       �                     *@        i       p                 ���"@������?
             1@       j       o                 ���!@z�G�z�?             $@       k       l                    �?      �?              @        ������������������������       �                     @        m       n                   �;@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        q       t                    ?@����X�?             @       r       s                   �<@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        w       �                    �?F��*���?           �z@        x       �                 �QD@��SK�?z            �g@       y       �                     @�BbΊ�?L             ]@        z       }                    �?     �?$             P@        {       |                     �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ~       �                    �?(;L]n�?"             N@              �                    :@��S�ۿ?             >@        �       �                   �5@"pc�
�?             &@        ������������������������       �                     @        �       �                   �3@�q�q�?             @       ������������������������       ����Q��?             @        ������������������������       �                     �?        ������������������������       �                     3@        ������������������������       �                     >@        �       �                    @��B����?(             J@       �       �                 ���4@�`���?%            �H@       �       �                    7@�!���?             A@        �       �                  �M$@�eP*L��?	             &@        ������������������������       �                      @        �       �                    �?�q�q�?             "@        ������������������������       �                     @        �       �                    �?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                   �;@��<b���?             7@        ������������������������       �                     "@        �       �                 ��.@X�Cc�?             ,@        �       �                   �<@���Q��?             @        ������������������������       �                      @        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                     @�<ݚ�?             "@       �       �                   �@@����X�?             @       �       �                    �?      �?             @        ������������������������       �                     �?        �       �                 ��1@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�r����?             .@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    @$�q-�?
             *@       ������������������������       �                     $@        �       �                    @�q�q�?             @        ������������������������       �                     �?        �       �                 ��T?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @`2U0*��?.            �R@       �       �                    �?�?�|�?-            �R@        ������������������������       �                    �A@        �       �                    �?�7��?            �C@       ������������������������       �                     ;@        �       �                    �?r�q��?             (@        ������������������������       �                      @        �       �                     @z�G�z�?             $@       �       �                    *@���Q��?             @        ������������������������       �                     �?        �       �                     �?      �?             @       �       �                   �>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �                           �?�j9:1w�?�            �m@        �       �                   �>@,ZYN(��?6            @T@        �       �                    �?V������?            �B@        �       �                  ��^@�t����?
             1@       �       �                    �?X�<ݚ�?             "@       �       �                   �:@      �?              @        ������������������������       �                      @        �       �                    =@�q�q�?             @       �       �                 �ܵ<@���Q��?             @        ������������������������       �                      @        �       �                 0��K@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �>@�z�G��?             4@        �       �                   �<@���Q��?             $@       �       �                   �;@և���X�?             @        ������������������������       �                     �?        �       �                 `fF<@      �?             @       �       �                 `fF:@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?z�G�z�?             $@       ������������������������       �                     @        �       �                    <@���Q��?             @       �       �                    7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                   �B@d�
��?             F@        �       �                    �?r�q��?             @       �       �                    �?�q�q�?             @        ������������������������       �                     �?        �       �                 03�P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �                          �?D�n�3�?             C@       �                          �?b�2�tk�?             B@       �       �                    �?*;L]n�?             >@        �       �                 @�pX@���Q��?             @       �       �                    �?      �?             @       �       �                 �̬L@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �                          �?���Q��?             9@       �       �                   �J@\X��t�?             7@       �       �                   �G@���Q��?	             .@       �       �                   �E@�q�q�?             "@        ������������������������       �                     �?        �       �                 `f�;@      �?              @       �       �                    G@�q�q�?             @       ������������������������       ����Q��?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                 `fF<@      �?              @       ������������������������       �                     @        �                        03wD@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @                                �K@r�q��?             @       ������������������������       �                     @                              `f�R@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        	                      ��&@Tݭg_�?b            �c@        
                      ��%@�q�q�?             (@                                 @�z�G��?             $@                               �5@�q�q�?             "@                                �1@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @                                 $@r�q��?[             b@                                  @X�<ݚ�?             ;@        ������������������������       �                     "@                              ��A>@r�q��?             2@        ������������������������       �                     "@                                 @�q�q�?             "@                                �?և���X�?             @        ������������������������       �                     @                                 @      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @                                 �9@��-�=��?I            @]@        ������������������������       �                     >@        !      6                   �?\-��p�?7            �U@        "      -                    @RB)��.�?            �E@       #      ,                ���,@�J�4�?             9@       $      +                  �D@      �?
             0@       %      &                  �;@���Q��?             $@        ������������������������       �                     �?        '      (                   �?X�<ݚ�?             "@        ������������������������       �                     �?        )      *                   @@      �?              @        ������������������������       �                     �?        ������������������������       �և���X�?             @        ������������������������       �                     @        ������������������������       �                     "@        .      5                   �?�E��ӭ�?             2@       /      0                   ;@�t����?             1@        ������������������������       �                     @        1      2                �T)D@؇���X�?
             ,@       ������������������������       �                     $@        3      4                   >@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     �?        7      B                  @@@t��ճC�?             F@       8      9                 �v6@�����H�?             ;@        ������������������������       �                     &@        :      A                   @     ��?             0@       ;      @                   �?�z�G��?             $@       <      =                039@�<ݚ�?             "@        ������������������������       �                     @        >      ?                  �?@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             1@        �t�bh�h*h-K ��h/��R�(KMCKK��h]�B0       �{@     �p@      m@     �I@      =@      >@       @      0@       @              @      0@      @      0@      @      @              @      @               @      *@               @       @      &@              @       @       @      �?              �?       @              �?      �?      @      �?      @              �?      �?              5@      ,@              @      5@       @      5@      @      *@      @      *@      @      @              "@      @      @      @      @       @      @       @       @              �?       @              �?      �?      �?      �?                      �?      @                       @      @                      �?       @                      @     �i@      5@     @f@      .@      a@      .@     @T@      (@      T@      $@      <@              J@      $@      $@              E@      $@       @      @               @       @      �?      �?              �?      �?      �?                      �?      D@      @      C@      @      "@              =@      @      <@      @      .@      �?      *@      �?      @      �?      �?              @      �?      @               @              *@      @      $@      @       @       @       @      �?              �?       @      �?      @              �?      �?      �?                      �?       @       @               @       @              �?       @      �?                       @     �K@      @              �?     �K@       @              �?     �K@      �?      7@              @@      �?      ?@      �?      ?@                      �?      �?              E@              :@      @      :@      @      *@              *@      @       @       @      @       @      @              @       @               @      @               @              @       @       @       @       @                       @      @                       @      j@     `k@     �@@     �c@      >@     �U@      @     �N@      �?      @      �?                      @       @      M@       @      <@       @      "@              @       @      @       @      @              �?              3@              >@      ;@      9@      8@      9@      &@      7@      @      @               @      @      @      @               @      @              @       @              @      2@              "@      @      "@      @       @       @              �?       @               @      �?               @      @       @      @       @       @              �?       @      �?              �?       @                      @               @      *@       @      �?      �?              �?      �?              (@      �?      $@               @      �?      �?              �?      �?      �?                      �?      @              @      R@       @      R@             �A@       @     �B@              ;@       @      $@               @       @       @       @      @      �?              �?      @      �?      �?      �?                      �?               @              @      �?              f@     �N@     �H@      @@      :@      &@      (@      @      @      @      @      @               @      @       @      @       @       @              �?       @               @      �?              �?                      �?       @              ,@      @      @      @      @      @              �?      @      @      @      �?      �?               @      �?               @      @               @       @      @              @       @      �?       @      �?                       @       @              7@      5@      �?      @      �?       @              �?      �?      �?              �?      �?                      @      6@      0@      6@      ,@      1@      *@       @      @      �?      @      �?      �?              �?      �?                       @      �?              .@      $@      *@      $@      @      "@      @      @              �?      @       @      @       @      @       @      �?               @                      @      @      �?      @               @      �?              �?       @               @              @      �?      @               @      �?       @                      �?               @     �_@      =@      @      @      @      @      @      @      �?      @      �?                      @      @              �?                       @      ^@      8@      .@      (@              "@      .@      @      "@              @      @      @      @      @              �?      @              @      �?               @             @Z@      (@      >@             �R@      (@      A@      "@      5@      @      (@      @      @      @      �?              @      @              �?      @      @      �?              @      @      @              "@              *@      @      (@      @              @      (@       @      $@               @       @       @      �?              �?      �?             �D@      @      8@      @      &@              *@      @      @      @      @       @      @               @       @       @                       @              �?      @              1@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ��(.hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM?huh*h-K ��h/��R�(KM?��h|�B�O         �                     @��"{��?�           @�@               _                    �?���Q��?�            `s@              8                     �?�85�r��?            �i@              5                    �?��̀�R�?C            �[@              $                   @F@<W#.m��?@            @Z@                                  �?z�7�Z�?/            @R@        ������������������������       �                    �A@               #                   @D@�����?             C@       	                          �<@V������?            �B@       
                           �?      �?             8@                                   �?؇���X�?             @                                  9@      �?             @        ������������������������       �                     �?                                03SA@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                `fF:@��.k���?	             1@        ������������������������       �                     @                                  �>@�q�q�?             (@        ������������������������       �                     @                                  �A@z�G�z�?             @        ������������������������       �                     @                                  `E@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               "                    �?8�Z$���?
             *@                                ��>@���Q��?             @        ������������������������       �                      @               !                    �?�q�q�?             @                                  �A@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        %       2                    �?      �?             @@       &       1                   �L@�û��|�?             7@       '       .                 03[=@�z�G��?             4@       (       )                    �?r�q��?             (@        ������������������������       �                      @        *       +                 ��:@z�G�z�?             $@        ������������������������       �                     �?        ,       -                   �J@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        /       0                   �@@      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        3       4                  DT@�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        6       7                    6@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        9       P                   @A@ާb�y��?<            �W@       :       O                    ?@և���X�?%             L@       ;       @                    �?
;&����?             G@        <       =                    �?և���X�?             @        ������������������������       �                     @        >       ?                 `��,@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        A       B                    @��
ц��?            �C@        ������������������������       �                     @        C       N                    �?��
P��?            �A@       D       E                    �?*;L]n�?             >@        ������������������������       �                     (@        F       G                    ;@�X�<ݺ?             2@       ������������������������       �                     "@        H       M                    �?�����H�?             "@       I       J                   �'@      �?              @        ������������������������       �                     @        K       L                    =@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        Q       ^                    �?�(�Tw��?            �C@       R       S                    �?<ݚ)�?             B@        ������������������������       �                     "@        T       U                    �?�>����?             ;@        ������������������������       �                     �?        V       [                   @N@$�q-�?             :@       W       Z                   @F@ �q�q�?             8@        X       Y                   @D@�C��2(�?             &@       ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                     *@        \       ]                   �P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        `       i                    �?���N8�?D            @Z@        a       h                    �? �.�?Ƞ?"             N@       b       g                    �?г�wY;�?             A@       c       f                   �6@      �?             @@        d       e                 ��m1@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     =@        ������������������������       �                      @        ������������������������       �                     :@        j       k                    +@��S���?"            �F@        ������������������������       �                     @        l       �                     �?p�ݯ��?             C@       m       �                    @� �	��?             9@       n       �                    �?�q�q�?             8@       o       �                    �?��Q��?             4@       p       q                   �;@p�ݯ��?             3@        ������������������������       �                     @        r                          �K@��S���?             .@       s       x                    �?��
ц��?
             *@        t       u                    C@�q�q�?             @        ������������������������       �                     �?        v       w                 @�pX@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        y       ~                 03�M@և���X�?             @       z       {                 �K@z�G�z�?             @        ������������������������       �                      @        |       }                 ��9L@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?      �?             @        ������������������������       �                      @        �       �                 `f�h@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        
             *@        �       �                    �?��5Е��?             y@        �       �                    >@ާb�y��?=            �W@       �       �                    @      �?8            �U@        ������������������������       �                     @        �       �                    @�W����?5            �T@       �       �                    �?z�G���?3             T@        �       �                 ��.@�E��ӭ�?             B@       �       �                   �-@��}*_��?             ;@        ������������������������       �                     �?        �       �                  S5&@$��m��?             :@       �       �                    �?���!pc�?             6@       �       �                    �?���N8�?
             5@        ������������������������       �                     @        �       �                   �8@     ��?             0@        ������������������������       �                      @        �       �                 ���@d}h���?             ,@        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                     �?        �       �                   �<@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        �       �                    �?v�X��?             F@       �       �                    �?$��m��?             :@       �       �                    �?���!pc�?             6@       �       �                    ;@z�G�z�?             .@        �       �                 xF*@      �?             @       �       �                 ���@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     &@        �       �                    �?և���X�?             @       �       �                    3@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �1@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                  ��@�<ݚ�?             2@        ������������������������       �                     @        �       �                 03�7@�	j*D�?	             *@       �       �                   �<@���|���?             &@       �       �                    �?�z�G��?             $@       �       �                    �?�<ݚ�?             "@       �       �                 ��(@      �?              @       ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     "@        �       �                    �?��Ji�?�            0s@        �       �                    �?7�A�0�?6             V@       �       �                    �?�;�vv��?,            @R@       �       �                   �;@X�<ݚ�?            �F@       �       �                    �?^������?            �A@       �       �                    9@\X��t�?             7@       �       �                 ���@�q�q�?
             .@        ������������������������       �                     @        �       �                  �#@�C��2(�?             &@       ������������������������       �                      @        �       �                 �[$@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?r�q��?             (@       �       �                    $@z�G�z�?             @        �       �                   �&@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ��l4@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                     @z�G�z�?             $@       �       �                   @"@      �?              @       ������������������������       �                     @        �       �                    I@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                   �B@��>4և�?             <@       �       �                   �>@�G��l��?             5@       �       �                   �.@����X�?             ,@        �       �                  S�$@�����H�?             "@        ������������������������       �                     @        �       �                    -@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    =@���Q��?             @       �       �                 pf�3@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    @��S�ۿ?
             .@       ������������������������       �                      @        �       �                    @؇���X�?             @        �       �                    @z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       8                �T�I@L��?�            `k@       �       7                   �?���H��?�            @j@       �       $                   �?(l58��?            �h@       �                         �3@�KM�]�?d             c@        �                          �2@z�G�z�?             9@       �       �                 ��Y @8�Z$���?             *@        �       �                    1@�q�q�?             @       �       �                 pf�@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                              �?�@      �?             (@        ������������������������       �                     @                              `�8"@�q�q�?             "@        ������������������������       �և���X�?             @        ������������������������       �                      @                              @3�@4Jı@�?U            �_@        ������������������������       �                      @                                �<@0{�v��?T            @_@       	                      ��L@��
���?0            �R@        
                      �?$@"pc�
�?	             &@                                ;@ףp=
�?             $@        ������������������������       �                     @                              pf�@z�G�z�?             @       ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �        '             P@              #                   �?�:pΈ��?$             I@                             �?�@8��8���?"             H@       ������������������������       �                     8@              "                  �G@�q�q�?             8@                               �>@�q�q�?             5@                                �=@�<ݚ�?             "@                             ���"@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @              !                @3�@�q�q�?	             (@                               �A@r�q��?             @        ������������������������       �                     @                                 �D@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        %      6                   �?��k=.��?            �G@       &      5                   0@���"͏�?            �B@       '      0                   �?      �?             8@       (      )                   3@�q�q�?             .@        ������������������������       �                     @        *      +                   5@�eP*L��?             &@        ������������������������       �                     @        ,      -                  �7@؇���X�?             @        ������������������������       �                     @        .      /                  �9@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        1      2                ���"@X�<ݚ�?             "@        ������������������������       �                     @        3      4                  �5@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     *@        ������������������������       �                     $@        ������������������������       �                     &@        9      >                p�O@�q�q�?             "@       :      =                   >@      �?              @       ;      <                   ;@���Q��?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     �?        �t�bh�h*h-K ��h/��R�(KM?KK��h]�B�       �y@     �r@      _@     @g@     �X@     �Z@     �G@     �O@      G@     �M@      :@     �G@             �A@      :@      (@      :@      &@      .@      "@      @      �?      @      �?      �?               @      �?              �?       @              @              "@       @      @              @       @              @      @      �?      @              �?      �?              �?      �?              &@       @      @       @       @              �?       @      �?      �?              �?      �?                      �?       @                      �?      4@      (@      ,@      "@      ,@      @      $@       @       @               @       @      �?              @       @               @      @              @      @              @      @                      @      @      @      @                      @      �?      @              @      �?              J@     �E@      8@      @@      8@      6@      @      @              @      @      �?              �?      @              5@      2@      @              1@      2@      1@      *@              (@      1@      �?      "@               @      �?      @      �?      @              @      �?              �?      @              �?                      @              $@      <@      &@      9@      &@              "@      9@       @      �?              8@       @      7@      �?      $@      �?       @               @      �?      *@              �?      �?              �?      �?              @              9@      T@      �?     �M@      �?     �@@      �?      ?@      �?       @               @      �?                      =@               @              :@      8@      5@              @      8@      ,@      &@      ,@      $@      ,@      @      *@      @      (@              @      @       @      @      @      @       @      �?              @       @               @      @              @      @      �?      @               @      �?       @      �?                       @       @                       @              �?      @      �?       @              �?      �?              �?      �?              �?              *@             0r@     �[@      J@     �E@     �E@     �E@              @     �E@     �C@     �D@     �C@      $@      :@      $@      1@      �?              "@      1@      @      0@      @      0@              @      @      &@       @              @      &@      @                      &@      �?              @      �?      @                      �?              "@      ?@      *@      1@      "@      0@      @      (@      @      �?      @      �?      �?              �?      �?                       @      &@              @      @      @      @              @      @              �?              �?      @      �?                      @      ,@      @      @              "@      @      @      @      @      @      @       @      @       @      @       @       @              �?                      �?              �?       @               @              "@             �m@      Q@     �I@     �B@     �B@      B@      4@      9@      (@      7@      $@      *@      $@      @              @      $@      �?       @               @      �?              �?       @                       @       @      $@      �?      @      �?      �?      �?                      �?              @      �?      @              @      �?               @       @      @       @      @              �?       @      �?                       @       @              1@      &@      $@      &@      $@      @       @      �?      @              @      �?              �?      @               @      @      �?      @              @      �?              �?                      @      @              ,@      �?       @              @      �?      @      �?      @                      �?       @             �g@      ?@      g@      9@     �e@      9@      a@      0@      4@      @      &@       @      @       @      @       @      @                       @      �?              @              "@      @      @              @      @      @      @       @              ]@      &@               @      ]@      "@     @R@       @      "@       @      "@      �?      @              @      �?      @              �?      �?              �?      P@             �E@      @     �D@      @      8@              1@      @      ,@      @      @       @      @       @      @                       @      @              @      @      �?      @              @      �?       @      �?      �?              �?      @              @               @              C@      "@      <@      "@      .@      "@      $@      @      @              @      @              @      @      �?      @              @      �?              �?      @              @      @      @               @      @              @       @              *@              $@              &@              @      @       @      @       @      @               @       @      �?              @      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJx�+hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM)huh*h-K ��h/��R�(KM)��h|�B@J         d                    �?z��Y�)�?�           @�@               ]                    @�]N���?�            @k@              "                  �#@.����?�             i@                                ���@�>$�*��?            �D@                                   1@���!pc�?
             &@        ������������������������       �                      @                                �Y�@�q�q�?             "@        ������������������������       �                      @        	       
                    9@؇���X�?             @        ������������������������       �                     @                                   �?      �?             @        ������������������������       �                     �?                                ���@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @               !                    K@�q�q�?             >@                                 �9@����X�?             <@                                   �?     ��?	             0@                               ���@@4և���?             ,@        ������������������������       �                      @                                   �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @                                   �?�q�q�?
             (@                                �&B@�q�q�?             @       ������������������������       ����Q��?             @        ������������������������       �                     �?                                   �@r�q��?             @                                  �A@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        #       \                    @��(\���?g             d@       $       M                 0#
9@
����?c             c@        %       0                     @z�z�7��?1            @R@       &       '                    �?Du9iH��?            �E@        ������������������������       �                     @        (       /                    �?�8��8��?             B@       )       .                    �?��2(&�?             6@       *       +                 `f�)@P���Q�?             4@        ������������������������       �                     @        ,       -                    :@@4և���?             ,@        ������������������������       ��q�q�?             @        ������������������������       �        
             &@        ������������������������       �                      @        ������������������������       �                     ,@        1       J                    �?�q�q�?             >@       2       =                    �?��X��?             <@        3       <                 ��l4@�z�G��?	             $@       4       ;                    �?�<ݚ�?             "@       5       :                 ���*@�q�q�?             @       6       9                    $@z�G�z�?             @        7       8                   �&@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        >       I                   �@@�q�q�?             2@       ?       @                    �?և���X�?	             ,@        ������������������������       �                     @        A       H                 ��1@�q�q�?             "@       B       C                    9@      �?             @        ������������������������       �                      @        D       E                   �.@      �?             @        ������������������������       �                      @        F       G                    ;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        K       L                  �2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        N       Y                    �?x�G�z�?2             T@       O       P                    �? ���J��?0            �S@        ������������������������       �                     =@        Q       R                    �?@9G��?            �H@        ������������������������       �                     4@        S       X                     �? 	��p�?             =@       T       U                    �?�r����?
             .@       ������������������������       �                     &@        V       W                 ���`@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     ,@        Z       [                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ^       _                     @@�0�!��?             1@        ������������������������       �                      @        `       c                    @��S�ۿ?             .@        a       b                    �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        e       �                     �?��_	f�?4           �~@        f       }                   �>@(Q����?A            @Y@        g       x                   �J@j���� �?             A@       h       i                    �?d��0u��?             >@        ������������������������       �                     @        j       w                   @D@l��
I��?             ;@       k       r                   �<@���Q��?
             4@       l       m                   �;@r�q��?             (@        ������������������������       �                      @        n       o                 �̌*@z�G�z�?             $@        ������������������������       �                     �?        p       q                 `fF<@�����H�?             "@        ������������������������       �      �?             @        ������������������������       �                     @        s       t                    A@      �?              @        ������������������������       �                     @        u       v                   �B@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        y       z                 `fF<@      �?             @        ������������������������       �                      @        {       |                   �P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ~       �                    �?.��<�?+            �P@              �                    �?���y4F�?%            �L@       �       �                   �A@     ��?             @@       �       �                    �?�E��ӭ�?             2@        �       �                    �?և���X�?             @       �       �                 0c@z�G�z�?             @        ������������������������       �                      @        �       �                   �?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                 ��yC@�C��2(�?             &@        �       �                   �@@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     ,@        �       �                 ��^@ �o_��?             9@       �       �                    D@      �?             8@        �       �                 �D�J@      �?              @        ������������������������       �                      @        �       �                    �?�q�q�?             @        �       �                 8�T@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �@@      �?             @        ������������������������       �                      @        �       �                 03U@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?      �?             0@        �       �                   �K@���Q��?             @       �       �                 @�pX@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     �?        �       �                    �?      �?             $@        ������������������������       �                     �?        �       �                     @X�<ݚ�?             "@       �       �                 ���i@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �G�?��w"��?�            �x@        ������������������������       �                     @        �                       ��T?@�cLN�)�?�            Px@       �                       �&@�I
��#�?�            �v@       �       
                �%@��d��?�            �o@       �       �                     @\�J��?�            @o@        �       �                   �5@�����?             5@        �       �                   �1@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        
             2@        �       �                 �?�@�H`}��?�            �l@       �       �                   �;@,I�e���?W            �b@        �       �                    �?     ��?#             P@       �       �                   �:@��[�8��?            �I@       �       �                 �Y�@r�q��?             H@        �       �                   �3@      �?
             0@        ������������������������       �                     @        �       �                    �?�n_Y�K�?             *@        �       �                 ��y@���Q��?             @        ������������������������       �                     �?        �       �                 ���@      �?             @        ������������������������       �                     �?        �       �                    5@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 �&b@      �?              @       �       �                 @33@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @@        ������������������������       �                     @        �       �                   �7@8�Z$���?             *@       ������������������������       �                     &@        ������������������������       �                      @        �       �                    �?`��F:u�?4            �U@        �       �                   @<@�C��2(�?             6@       �       �                 ���@8�Z$���?             *@        ������������������������       �                     @        �       �                   @@�q�q�?             @       ������������������������       �      �?             @        ������������������������       �                      @        ������������������������       �                     "@        �       �                   �<@��ɉ�?&            @P@        ������������������������       �                     A@        �       �                   �=@`Jj��?             ?@        ������������������������       �                     �?        �       �                    �?(;L]n�?             >@        ������������������������       �                     @        �       �                 �&B@ �q�q�?             8@       ������������������������       �                     4@        �       �                   �@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �:@����?4            �S@        �       �                    �?��� ��?             ?@       �       �                 ��Y @�r����?             >@       �       �                 @3�@������?             1@        ������������������������       �                      @        �       �                   �3@������?	             .@        �       �                   �1@�q�q�?             @        ������������������������       �                      @        ������������������������       �      �?             @        ������������������������       �                     "@        ������������������������       �        
             *@        ������������������������       �                     �?        �       	                   �?(���@��?            �G@       �       �                 @3�@�I� �?             G@        �       �                   �?@��S���?             .@        ������������������������       �                      @        �       �                   �D@��
ц��?             *@       �       �                   @A@���|���?             &@        ������������������������       �և���X�?             @        �       �                    C@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                      @        �       �                    �?��a�n`�?             ?@        ������������������������       �                     �?        �       �                   �;@�������?             >@        ������������������������       �                     �?        �                       ��) @V�a�� �?             =@       �       �                    ?@P���Q�?             4@       ������������������������       �        	             .@                                 �@@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @                                 ?@X�<ݚ�?             "@                              `��!@r�q��?             @        ������������������������       �                     @                              ���"@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @                                 �?�/�z{�?H            @\@                               �*@����D��?8            @W@                                �>@      �?             @@                                �?؇���X�?
             ,@                               �;@8�Z$���?	             *@       ������������������������       �                     &@        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     2@        ������������������������       �        &            �N@                              03{3@ףp=
�?             4@                              `ff/@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     .@              (                  �?@�q�q�?             8@             !                   �?��s����?             5@                              �DpB@ףp=
�?	             $@                                 +@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        "      #                   �?���!pc�?             &@        ������������������������       �                     �?        $      '                   @�z�G��?             $@        %      &                pf�C@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �t�b��     h�h*h-K ��h/��R�(KM)KK��h]�B�       �|@     @o@      N@     �c@      G@     `c@      7@      2@      @       @               @      @      @       @              �?      @              @      �?      @              �?      �?       @      �?                       @      4@      $@      4@       @      *@      @      *@      �?       @              @      �?              �?      @                       @      @      @       @      @       @      @              �?      @      �?      �?      �?              �?      �?              @                       @      7@      a@      0@      a@      *@      N@      @      D@              @      @     �@@      @      3@      �?      3@              @      �?      *@      �?       @              &@       @                      ,@      $@      4@      "@      3@      @      @       @      @       @      @      �?      @      �?      �?      �?                      �?              @      �?                      @      �?              @      (@      @       @              @      @      @      @      @               @      @      �?       @              �?      �?      �?                      �?      @                      @      �?      �?      �?                      �?      @     @S@       @      S@              =@       @     �G@              4@       @      ;@       @      *@              &@       @       @               @       @                      ,@      �?      �?              �?      �?              @              ,@      @               @      ,@      �?      @      �?              �?      @               @              y@      W@      P@     �B@      ,@      4@      &@      3@      @               @      3@       @      (@       @      $@               @       @       @      �?              �?       @      �?      @              @      @       @      @              @       @               @      @                      @      @      �?       @              �?      �?      �?                      �?      I@      1@     �F@      (@      ;@      @      *@      @      @      @      �?      @               @      �?       @      �?                       @       @              $@      �?      @      �?      @                      �?      @              ,@              2@      @      2@      @      @      @       @               @      @      �?      �?              �?      �?              �?      @               @      �?      �?      �?                      �?      ,@       @      @       @      @      �?              �?      @                      �?      &@                      �?      @      @              �?      @      @      �?      @              @      �?              @              u@     �K@              @      u@     �I@     t@      F@     �j@      D@     �j@      C@      3@       @      �?       @      �?                       @      2@              h@      B@     �`@      1@     �I@      *@      D@      &@      D@       @       @       @      @              @       @       @      @      �?              �?      @              �?      �?       @               @      �?              @      @      @       @               @      @                      @      @@                      @      &@       @      &@                       @     �T@      @      4@       @      &@       @      @              @       @       @       @       @              "@             �O@       @      A@              =@       @              �?      =@      �?      @              7@      �?      4@              @      �?              �?      @             �M@      3@      ;@      @      :@      @      *@      @       @              &@      @       @      @               @       @       @      "@              *@              �?              @@      .@      ?@      .@      @       @               @      @      @      @      @      @      @      @      �?      �?               @      �?               @      8@      @      �?              7@      @              �?      7@      @      3@      �?      .@              @      �?              �?      @              @      @      �?      @              @      �?       @      �?                       @      @              �?                       @     @[@      @     �V@       @      >@       @      (@       @      &@       @      &@                       @      �?              2@             �N@              2@       @      @       @      @                       @      .@              1@      @      1@      @      "@      �?      �?      �?              �?      �?               @               @      @      �?              @      @       @      @              @       @              @                      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJH�SshG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B�B         `                    �?b�`�6��?�           @�@                                `f�$@`�B7��?�             p@                                   �?և���X�?"            �H@        ������������������������       �                     @                                   @F�����?            �F@                                  A@8�$�>�?            �E@                                 �>@\�Uo��?             C@                                  �?*O���?             B@       	                        pF @     ��?             @@       
                           @���Q��?             4@        ������������������������       �                      @                                 s�@�q�q�?             2@        ������������������������       �                     @                                   �?      �?
             (@                                 �5@�q�q�?             "@        ������������������������       �                     �?                                   �?      �?              @                               �&B@r�q��?             @       ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @                                   3@�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @               I                    �?J�B�9��?�             j@              B                 м�9@��V���?^            �c@               A                    @ڤ���?1            @T@       !       ,                 �B,@��n�?.            �R@        "       +                     @P�Lt�<�?             C@       #       *                    �?(;L]n�?             >@       $       %                 `f�)@XB���?             =@        ������������������������       �                     &@        &       )                   �*@�X�<ݺ?             2@       '       (                    :@      �?	             0@        ������������������������       �                     �?        ������������������������       �                     .@        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        -       @                    �?^H���+�?            �B@       .       /                    .@�P�*�?             ?@        ������������������������       �                     @        0       9                    �? �o_��?             9@       1       2                    �?և���X�?	             ,@        ������������������������       �                     @        3       6                   �;@�eP*L��?             &@        4       5                 @3�/@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        7       8                 03�1@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        :       ?                   �>@�C��2(�?             &@        ;       <                    �?z�G�z�?             @        ������������������������       �                     @        =       >                     @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        C       D                   �H@P�Lt�<�?-             S@       ������������������������       �        %             P@        E       H                   @I@r�q��?             (@        F       G                     �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        J       W                 03�;@��WV��?$             J@        K       V                    @�㙢�c�?             7@       L       S                 ��97@��2(&�?             6@       M       R                    �?@4և���?	             ,@        N       Q                   �<@      �?             @       O       P                 `�@1@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        T       U                 039@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        X       _                     @J�8���?             =@       Y       Z                    �?����X�?             ,@        ������������������������       �                      @        [       ^                     @�q�q�?	             (@       \       ]                 ���`@���Q��?             $@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        
             .@        a       j                    @�.U֪E�?-           `|@        b       g                    �?      �?             8@       c       d                 ���3@j���� �?             1@        ������������������������       �                     @        e       f                    @���|���?             &@        ������������������������       �                     @        ������������������������       �                     @        h       i                    @����X�?             @       ������������������������       �                     @        ������������������������       �                      @        k       �                 ��D:@�g��?           �z@       l       }                     @@[�f�?�            �s@        m       n                     �? �q�q�?5             R@        ������������������������       �                     @        o       |                   �*@P�2E��?0            @P@       p       q                    �?@4և���?             E@        ������������������������       �                     �?        r       s                 `fF)@��p\�?            �D@        ������������������������       �                     3@        t       u                   �;@��2(&�?             6@        ������������������������       �                     $@        v       w                    =@      �?             (@        ������������������������       �                      @        x       {                   @B@ףp=
�?             $@       y       z                    @@      �?             @        ������������������������       �                      @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     7@        ~       �                    �?l���u�?�            `n@               �                    ;@8�Z$���?            �C@        �       �                 �&2.@�q�q�?             (@       �       �                    �?r�q��?             @       �       �                 ���@z�G�z�?             @        ������������������������       �                      @        �       �                 H�%@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?�q�q�?             @       �       �                   �2@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   @<@ 7���B�?             ;@       �       �                 ���@�IєX�?             1@        ������������������������       �                     @        �       �                   @@ףp=
�?             $@       ������������������������       �؇���X�?             @        ������������������������       �                     @        ������������������������       �                     $@        �       �                    �?`�H�/��?}            �i@       �       �                   @C@��-�=��?u            `h@       �       �                   �;@l��\��?f            @e@        �       �                    �?��2(&�?(            �P@        ������������������������       �                     @        �       �                    �?���-T��?&             O@       �       �                   �:@X�;�^o�?"            �K@       �       �                   �8@@�E�x�?             �H@       ������������������������       �                     E@        �       �                   �9@؇���X�?             @        �       �                 @33@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �6@����X�?             @        �       �                   �2@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                 ��@0G���ջ?>             Z@        ������������������������       �                     <@        �       �                    �?�˹�m��?/             S@       �       �                   @@@���}<S�?+            @Q@       �       �                   �<@�KM�]�?%            �L@       �       �                    �?���.�6�?             G@        ������������������������       �                     @        �       �                 �?$@@4և���?             E@        ������������������������       �                      @        �       �                 ��) @�(\����?             D@       ������������������������       �                     <@        �       �                 pf� @�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        �       �                   �=@���!pc�?             &@        �       �                 �̌!@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                   �@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        ������������������������       �                     @        �       �                   �C@z�G�z�?             9@        ������������������������       �      �?             @        �       �                   @F@�����?             5@        �       �                 ��Y@����X�?             @        ������������������������       �                     @        �       �                 pf� @      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        	             ,@        ������������������������       �                     "@        �                          �?pi�hv#�?P            �\@       �       �                    �?PN���?B            @V@       �       �                 `f�B@�q�q�?,            �L@        �       �                    �?      �?             >@       �       �                 ���=@���>4��?             <@       �       �                 03k:@�q�q�?             .@        ������������������������       �                      @        �       �                    J@�θ�?             *@       �       �                   `G@      �?              @       �       �                    �?����X�?             @        ������������������������       �                      @        �       �                   �F@���Q��?             @       �       �                   @B@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �>@�θ�?             *@       ������������������������       �                      @        �       �                   �@@���Q��?             @        ������������������������       �                     �?        �       �                   @B@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?PN��T'�?             ;@       �       �                   �?@z�G�z�?             4@       �       �                    �?�r����?             .@        ������������������������       �                     @        �       �                      @z�G�z�?	             $@       ������������������������       �                     @        �       �                    ;@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        �       �                   �A@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �                        D�\@     ��?             @@       �       �                 03U@V�a�� �?             =@       �       �                    +@�J�4�?             9@        ������������������������       �                     �?        �       �                     �?      �?             8@        �       �                    �?�θ�?             *@       �       �                   @K@ףp=
�?             $@        �       �                    7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                  x�N@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        �                          �?      �?             @                                 F@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                 �? ��WV�?             :@        ������������������������       �                      @                              ���Y@ �q�q�?             8@       ������������������������       �        
             6@        	      
                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �t�bh�h*h-K ��h/��R�(KMKK��h]�B�       `|@      p@     @R@      g@      <@      5@              @      <@      1@      <@      .@      7@      .@      7@      *@      3@      *@       @      (@       @              @      (@              @      @      @      @      @              �?      @      @      �?      @      �?       @              @       @              @              &@      �?              �?      &@              @                       @      @                       @     �F@     �d@      6@     �`@      4@     �N@      ,@     �N@      �?     �B@      �?      =@      �?      <@              &@      �?      1@      �?      .@      �?                      .@               @              �?               @      *@      8@      *@      2@      @              @      2@      @       @              @      @      @      @      �?              �?      @               @      @              @       @              �?      $@      �?      @              @      �?      �?              �?      �?                      @              @      @               @     �R@              P@       @      $@       @       @       @                       @               @      7@      =@      @      3@      @      3@      �?      *@      �?      @      �?      �?      �?                      �?               @              $@       @      @       @                      @      �?              3@      $@      @      $@               @      @       @      @      @              @      @                       @      .@             �w@     @R@      "@      .@      @      $@              @      @      @              @      @               @      @              @       @             @w@      M@     �q@      =@     @Q@      @      @              O@      @     �C@      @      �?              C@      @      3@              3@      @      $@              "@      @               @      "@      �?      @      �?       @              �?      �?      @              7@              k@      :@     �@@      @      @      @      @      �?      @      �?       @               @      �?              �?       @              �?               @      @       @      @       @                      @              �?      :@      �?      0@      �?      @              "@      �?      @      �?      @              $@              g@      4@     �e@      4@     `c@      .@     �L@      "@      @             �J@      "@      H@      @      H@      �?      E@              @      �?      @      �?              �?      @              @                      @      @       @       @       @       @                       @      @             �X@      @      <@             �Q@      @     �O@      @     �I@      @     �E@      @      @             �C@      @               @     �C@      �?      <@              &@      �?              �?      &@               @      @      @       @      @                       @      @      �?              �?      @              (@              @              4@      @      �?      @      3@       @      @       @      @               @       @               @       @              ,@              "@             �U@      =@     �N@      <@      C@      3@      .@      .@      *@      .@      $@      @               @      $@      @      @      @      @       @       @              @       @      �?       @      �?      �?              �?       @                      �?      @              @      $@               @      @       @      �?               @       @               @       @               @              7@      @      0@      @      *@       @      @               @       @      @               @       @              �?       @      �?      @       @               @      @              @              7@      "@      7@      @      5@      @              �?      5@      @      $@      @      "@      �?       @      �?       @                      �?      @              �?       @               @      �?              &@               @       @      �?       @               @      �?              �?                      @      9@      �?       @              7@      �?      6@              �?      �?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�8�hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMAhuh*h-K ��h/��R�(KMA��h|�B@P         x                  �#@�U��h��?�           @�@               /                    �?h��Q(�?�            �p@                                P��@h�n��?2            @U@                                ��Y@������?             A@        ������������������������       �                     @                                   5@�c�Α�?             =@        ������������������������       �                      @                                   �?�<ݚ�?             ;@        	       
                    �?      �?              @       ������������������������       �                     @        ������������������������       �                     @                                   �?�}�+r��?             3@                               ���@�IєX�?             1@                                 �7@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     @        ������������������������       �                      @                                   �?j���� �?            �I@                                �� @      �?              @                                  ?@����X�?             @                                 �<@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?               .                    �?�+��<��?            �E@              '                    �?D^��#��?            �D@                                  �2@R���Q�?             4@        ������������������������       �                     @               &                 �&B@@�0�!��?
             1@               !                  s�@�θ�?             *@        ������������������������       �                      @        "       #                   �5@���!pc�?             &@        ������������������������       �                     �?        $       %                    9@z�G�z�?             $@        ������������������������       �                     �?        ������������������������       ��<ݚ�?             "@        ������������������������       �                     @        (       )                  ��@�����?             5@        ������������������������       �                     @        *       -                 ��(@      �?             0@       +       ,                   �=@؇���X�?             ,@       ������������������������       ��<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        0       C                    �?f>�cQ�?u            �f@        1       2                    3@�q�q�?             5@        ������������������������       �                     �?        3       4                 ���@�z�G��?             4@        ������������������������       �                      @        5       B                    �?�<ݚ�?             2@       6       A                    K@������?             .@       7       @                  SE"@d}h���?
             ,@       8       ?                 ��� @�z�G��?             $@       9       :                   �6@�<ݚ�?             "@        ������������������������       �                     �?        ;       >                    ;@      �?              @        <       =                   �9@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        D       w                   �C@�$�����?e            @d@       E       r                    �?��8���?Y            �a@       F       G                     @�LQ�1	�?T            @a@        ������������������������       �                     "@        H       q                   @C@(L���?O             `@       I       \                 �?�@ ��P0�?N            �_@       J       [                   �;@�#-���?-            �Q@       K       N                 ��@�S����?             C@        L       M                    7@      �?             @        ������������������������       �                      @        ������������������������       �                      @        O       Z                   �:@�t����?             A@       P       Y                 �1@�C��2(�?            �@@       Q       R                   �4@؇���X�?             5@        ������������������������       �                      @        S       T                   �5@�θ�?
             *@        ������������������������       �                      @        U       V                    7@�C��2(�?	             &@        ������������������������       �                     @        W       X                   �8@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             (@        ������������������������       �                     �?        ������������������������       �                     @@        ]       j                   �<@�k�'7��?!            �L@       ^       e                   �3@��2(&�?             F@        _       d                   �2@�θ�?             *@       `       c                   �0@�����H�?             "@       a       b                 pFD!@r�q��?             @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �      �?             @        f       g                 ��) @��a�n`�?             ?@       ������������������������       �        
             1@        h       i                 pf� @d}h���?             ,@        ������������������������       �                     @        ������������������������       �                     &@        k       n                   �=@�	j*D�?             *@        l       m                 ���"@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        o       p                 @3�@z�G�z�?             $@        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                      @        s       v                    �?���Q��?             @       t       u                   �:@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     3@        y       �                    �?r�J���?            �{@        z       �                     @��3E��?|            @g@       {       �                    �?PF��t<�?U            �_@       |       }                     �?��F�D�?D            �X@       ������������������������       �        %             L@        ~       �                    �? �#�Ѵ�?            �E@              �                   �;@ 	��p�?             =@        �       �                   �6@�<ݚ�?             "@        ������������������������       �                     @        �       �                   �7@���Q��?             @       �       �                   �9@�q�q�?             @        ������������������������       �                     �?        �       �                   �/@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     4@        ������������������������       �                     ,@        �       �                    @@4և���?             <@       �       �                 ���`@�>����?             ;@       ������������������������       �                     4@        �       �                    �?����X�?             @       �       �                 Ъ�c@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�m����?'            �M@       �       �                    @v�2t5�?            �D@       �       �                    �?">�֕�?            �A@        �       �                    "@      �?              @        ������������������������       �                      @        �       �                    5@�q�q�?             @        ������������������������       �                     @        �       �                    :@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 `f7@������?             ;@       �       �                    �?z�G�z�?             9@        ������������������������       �                     @        �       �                   �D@�GN�z�?             6@       �       �                    =@��s����?             5@       �       �                   @.@      �?             0@       �       �                    �?���Q��?             $@       �       �                    $@����X�?             @        �       �                   �&@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 �[$@z�G�z�?             @        ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    -@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�E��ӭ�?             2@        ������������������������       �                      @        �       �                 pfv2@     ��?             0@        ������������������������       �                      @        �       �                    �?@4և���?
             ,@        ������������������������       �                     @        �       �                    @�C��2(�?             &@        �       �                 ��T?@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       .                 D0T@`�B7��?�             p@       �       �                    �?�1�d��?�             l@        �       �                 @Q,@�z�G��?             >@        ������������������������       �                     @        �       �                     �?���B���?             :@       �       �                   �;@      �?
             0@        ������������������������       �                      @        �       �                   �J@؇���X�?             ,@       �       �                    �?$�q-�?             *@       �       �                    ?@�C��2(�?             &@       ������������������������       �                     "@        �       �                    A@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                     @ףp=
�?	             $@        ������������������������       �                     @        �       �                    ;@r�q��?             @       �       �                 �0@�q�q�?             @        ������������������������       �                     �?        �       �                   �2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       -                `f�N@�U�u]�?~            `h@       �       &                �TL@      �?r             f@       �       �                     �?x���@O�?n             e@        �       �                    �?���Q��?            �F@       �       �                   �F@D�n�3�?             C@       �       �                   �@@\X��t�?             7@       �       �                   �>@�\��N��?             3@        �       �                   �<@z�G�z�?             $@       �       �                   �;@�����H�?             "@        ������������������������       �                     @        �       �                 `fF<@r�q��?             @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �=@�����H�?             "@       �       �                   �A@؇���X�?             @        ������������������������       �                     @        �       �                 ��yC@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    R@z�G�z�?	             .@       �       �                   @J@$�q-�?             *@        �       �                   �H@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                   @K@����X�?             @       �       �                  x#J@      �?             @        ������������������������       �                     �?        �       �                 `�iJ@�q�q�?             @        ������������������������       �                     �?        �       �                    7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                  �?�חF�P�?Q             _@                                 �?؇���X�?             ,@        ������������������������       �                     @                                 �?����X�?             @        ������������������������       �                      @        ������������������������       �                     @                                 !@�2����?I            �[@                                 �?�<ݚ�?             2@                               C@     ��?	             0@       	      
                ���3@@4և���?             ,@        ������������������������       �                     @                                  @؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @                                 @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?              %                   0@�nkK�?>             W@              $                `ff.@������?            �B@             #                    @�8��8��?             B@                                &@��a�n`�?             ?@                                �5@8�Z$���?             *@                                �1@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     "@                                �(@�X�<ݺ?             2@        ������������������������       �                     �?                                 C@�IєX�?             1@       ������������������������       �                     "@              "                  �*@      �?              @              !                  �F@؇���X�?             @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        #            �K@        '      ,                   �?؇���X�?             @       (      )                   ;@z�G�z�?             @        ������������������������       �                      @        *      +                   >@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     3@        /      >                03c@����e��?            �@@       0      =                   �?"pc�
�?             6@       1      <                   �?�q�q�?             (@       2      3                   �?���Q��?             $@        ������������������������       �                     �?        4      5                  �:@�q�q�?             "@        ������������������������       �                     @        6      ;                   �?      �?             @       7      8                  @C@���Q��?             @        ������������������������       �                     �?        9      :                @�pX@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        ?      @                @�:x@"pc�
�?             &@       ������������������������       �                     "@        ������������������������       �                      @        �t�bh�h*h-K ��h/��R�(KMAKK��h]�B       �z@     �q@     �j@      L@      L@      =@      :@       @      @              5@       @               @      5@      @      @      @              @      @              2@      �?      0@      �?      "@      �?              �?      "@              @               @              >@      5@      @       @      @       @       @       @       @                       @      @              �?              8@      3@      6@      3@      @      1@              @      @      ,@      @      $@               @      @       @      �?               @       @              �?       @      @              @      3@       @      @              ,@       @      (@       @      @       @      @               @               @             �c@      ;@      ,@      @              �?      ,@      @               @      ,@      @      &@      @      &@      @      @      @      @       @              �?      @      �?       @      �?       @                      �?      @                      �?      @                      �?      @             �a@      4@     �^@      4@      ^@      2@      "@             �[@      2@     �[@      0@      P@      @      @@      @       @       @       @                       @      >@      @      >@      @      2@      @       @              $@      @               @      $@      �?      @              @      �?              �?      @              (@                      �?      @@             �G@      $@      C@      @      $@      @       @      �?      @      �?      �?      �?      @              @               @       @      <@      @      1@              &@      @              @      &@              "@      @      �?       @      �?                       @       @       @       @       @      @                       @      @       @       @       @               @       @              �?              3@             `k@      l@      A@      c@      @     �^@       @     @X@              L@       @     �D@       @      ;@       @      @              @       @      @       @      �?      �?              �?      �?              �?      �?                       @              4@              ,@       @      :@       @      9@              4@       @      @       @      �?       @                      �?              @              �?      >@      =@      1@      8@      &@      8@      @      @               @      @       @      @              �?       @               @      �?              @      4@      @      4@              @      @      1@      @      1@      @      (@      @      @       @      @      �?      �?      �?                      �?      �?      @              @      �?      �?      �?                      �?       @      �?              �?       @                      @              @      �?               @              @              *@      @               @      *@      @               @      *@      �?      @              $@      �?       @      �?       @                      �?       @              g@     @R@     �e@     �J@      5@      "@              @      5@      @      (@      @               @      (@       @      (@      �?      $@      �?      "@              �?      �?              �?      �?               @                      �?      "@      �?      @              @      �?       @      �?      �?              �?      �?      �?                      �?      @             �b@      F@     �`@      F@     ``@      C@      ;@      2@      6@      0@      $@      *@      $@      "@       @       @      �?       @              @      �?      @      �?      �?              @      �?               @      �?      @      �?      @              @      �?              �?      @               @                      @      (@      @      (@      �?      @      �?      @                      �?       @                       @      @       @       @       @      �?              �?       @              �?      �?      �?      �?                      �?      @              Z@      4@      (@       @      @              @       @               @      @              W@      2@      @      ,@      @      *@      �?      *@              @      �?      @              @      �?               @              �?      �?              �?      �?              V@      @     �@@      @     �@@      @      <@      @      &@       @       @       @      �?              �?       @      "@              1@      �?      �?              0@      �?      "@              @      �?      @      �?       @      �?      @              �?              @                      �?     �K@              �?      @      �?      @               @      �?       @      �?                       @               @      3@              *@      4@      @      2@      @       @      @      @      �?              @      @              @      @      @       @      @      �?              �?      @              @      �?              �?                       @              $@      "@       @      "@                       @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJUehG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B�G         b                    �?l��n�?�           @�@                                    @\F~�1�?�            �n@                                   �?H�Swe�?P            @_@                                 �;@ ��Ou��?4            �S@                                  �7@؇���X�?             5@                                  �7@      �?             @        ������������������������       �                      @               	                    �?      �?             @        ������������������������       �                     �?        
                        ��m1@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     .@                                   �?���U�?$            �L@                                ��A@�r����?             .@        ������������������������       �                      @        ������������������������       �        
             *@        ������������������������       �                     E@                                   @`Ql�R�?            �G@        ������������������������       �                     �?        ������������������������       �                     G@               [                    @��S���?R             ^@              6                    �?���r
��?D            @X@               +                    �?�<ݚ�?            �F@              $                   �5@@�0�!��?             A@                                03�@�q�q�?             (@        ������������������������       �                      @                                   �?�z�G��?             $@                                ��%@      �?             @        ������������������������       �                     @        ������������������������       �                     �?                !                  s�@�q�q�?             @        ������������������������       �                      @        "       #                    2@      �?             @        ������������������������       �                      @        ������������������������       �                      @        %       &                    9@���7�?             6@        ������������������������       �                      @        '       *                    �?P���Q�?             4@        (       )                 H�%@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     1@        ,       -                    &@���|���?	             &@        ������������������������       �                     @        .       5                    @և���X�?             @       /       0                 03�-@�q�q�?             @        ������������������������       �                     @        1       4                  S�2@�q�q�?             @       2       3                   �<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        7       Z                    �?��
ц��?'             J@       8       O                 `f�%@�q�����?%             I@       9       :                 ���@     ��?             @@        ������������������������       �                     @        ;       J                 @3�"@>���Rp�?             =@       <       I                    �?�q�q�?             2@       =       D                   �;@�t����?             1@       >       A                 P�@X�<ݚ�?             "@        ?       @                    4@      �?             @        ������������������������       �                      @        ������������������������       �                      @        B       C                   �9@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        E       F                   �>@      �?              @       ������������������������       �                     @        G       H                    C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        K       L                 Ь�#@�C��2(�?             &@        ������������������������       �                     @        M       N                  �M$@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        P       Y                 `f68@�<ݚ�?             2@       Q       X                    �?      �?             0@       R       W                   @C@�q�q�?             @       S       T                 @3�/@z�G�z�?             @        ������������������������       �                      @        U       V                    ;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                      @        ������������������������       �                      @        \       ]                 pfv2@��<b���?             7@        ������������������������       �                      @        ^       a                    @؇���X�?             5@       _       `                 ��T?@d}h���?             ,@       ������������������������       �                     &@        ������������������������       �                     @        ������������������������       �                     @        c       �                 ���=@�5*S��?#           0}@       d       �                    �?hau��?�            �v@       e       �                   �<@H%u��?�            Pt@       f       �                   �5@�����?}            �h@        g       z                   �3@t/*�?             �G@       h       i                    �?ܷ��?��?             =@        ������������������������       �                     @        j       s                   �2@ȵHPS!�?             :@        k       l                     @@4և���?	             ,@        ������������������������       �                     @        m       r                    �?؇���X�?             @       n       q                   �0@z�G�z�?             @        o       p                 pf�@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        t       u                     @r�q��?	             (@        ������������������������       �      �?              @        v       w                 �?�@ףp=
�?             $@       ������������������������       �                     @        x       y                 `�8"@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        {       �                    �?�E��ӭ�?             2@       |                           �?������?             1@        }       ~                 �{@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 �1@؇���X�?
             ,@        �       �                  s@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �                     �?        �       �                   �8@�E�0�/�?]             c@        ������������������������       �                    �D@        �       �                    �?̹�"���?K            �[@        �       �                 @Q,@R���Q�?             4@       �       �                   @<@�z�G��?             $@       �       �                 ��%@�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        �       �                   �;@|)����??            �V@        �       �                 ��]@�+e�X�?             9@        �       �                   �:@X�<ݚ�?             "@       �       �                    �?�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �:@      �?             0@       ������������������������       �        	             *@        �       �                     @�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                 pf� @Pa�	�?-            �P@       �       �                    �?�nkK�?             G@        �       �                  s�@$�q-�?             *@        ������������������������       �                     @        �       �                    �?      �?              @       ������������������������       �z�G�z�?             @        ������������������������       �                     @        �       �                 ��) @Pa�	�?            �@@       ������������������������       �                     @@        ������������������������       �                     �?        ������������������������       �                     4@        �       �                     @��d��?L            �_@        �       �                 ��$:@�j��b�?!            �M@       �       �                    �?�7��?            �C@       �       �                    �? >�֕�?            �A@        ������������������������       �                      @        �       �                   �'@�FVQ&�?            �@@        ������������������������       �                     ,@        �       �                     �?�KM�]�?             3@        ������������������������       �                     �?        �       �                   @B@�����H�?
             2@        �       �                    @@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     *@        ������������������������       �                     @        �       �                 03k:@z�G�z�?             4@        ������������������������       �                      @        �       �                    H@�����H�?
             2@        ������������������������       �                     "@        �       �                   �J@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?h��Q(�?+            �P@       �       �                 �&B@�<ݚ�?(            �O@        �       �                 ���@`2U0*��?             9@       ������������������������       �                     1@        �       �                    >@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   @@@P����?             C@        �       �                    �?X�Cc�?	             ,@        ������������������������       �                     �?        �       �                   �>@�n_Y�K�?             *@        �       �                   �=@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �?�@�<ݚ�?             "@        �       �                   �@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �?@؇���X�?             @        ������������������������       �                     @        �       �                 @3�@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        �       �                   @C@r�q��?             8@        ������������������������       �                     (@        �       �                   �F@�q�q�?             (@       �       �                 @3�@      �?              @       �       �                   �D@z�G�z�?             @       ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    :@D^��#��?            �D@       �       �                    �?     ��?             @@        ������������������������       �                     @        �       �                 ���#@���>4��?             <@        ������������������������       �                     @        �       �                    0@�LQ�1	�?             7@       �       �                     @      �?	             0@       ������������������������       �                     .@        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        �                          @n�ޢ
�?A            @Y@       �                          @�ҿf���?7            �T@       �       �                   �1@D^��#��?6            �T@        ������������������������       �                     @        �       �                    @@��Zy�?3            �S@        �       �                     �?d}h���?	             ,@       �       �                   @>@8�Z$���?             *@        �       �                   @K@r�q��?             @       �       �                   �<@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �J@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �                          >@     x�?*             P@        �                           @�n`���?             ?@       �                          �?�����?             5@       �                       �U�X@"pc�
�?             &@        �                          �?���Q��?             @       �       �                    �?      �?             @        ������������������������       �                     �?                                 �U@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@                                 ;@���Q��?             $@        ������������������������       �                     �?        ������������������������       ��q�q�?             "@        	                          @�'�=z��?            �@@       
                         �?��S���?             >@                                 �?�z�G��?             $@                                �?      �?              @        ������������������������       �                     @                              @�pX@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @                                �F@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                 �?��Q��?             4@        ������������������������       �                     @                                  �?��
ц��?             *@                                �?�z�G��?             $@                               @K@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             2@        �t�b�      h�h*h-K ��h/��R�(KMKK��h]�B�       {@     pq@      O@     �f@      @     �]@      @     @R@      @      2@      @      @               @      @      �?      �?               @      �?              �?       @                      .@       @     �K@       @      *@       @                      *@              E@      �?      G@      �?                      G@      L@      P@      C@     �M@      $@     �A@      @      <@      @      @       @              @      @      �?      @              @      �?               @      @               @       @       @               @       @              �?      5@               @      �?      3@      �?       @               @      �?                      1@      @      @              @      @      @      @       @      @              �?       @      �?      �?      �?                      �?              �?              �?      <@      8@      :@      8@      6@      $@              @      6@      @      (@      @      (@      @      @      @       @       @       @                       @      @       @      @                       @      @      �?      @              �?      �?              �?      �?                      �?      $@      �?      @              @      �?              �?      @              @      ,@       @      ,@       @      @      �?      @               @      �?       @      �?                       @      �?                      $@       @               @              2@      @               @      2@      @      &@      @      &@                      @      @             0w@      X@     @s@      M@     �q@     �C@     �f@      3@     �C@       @      :@      @      @              7@      @      *@      �?      @              @      �?      @      �?       @      �?       @                      �?       @               @              $@       @      �?      �?      "@      �?      @              @      �?              �?      @              *@      @      *@      @      �?       @      �?                       @      (@       @       @       @       @                       @      $@                      �?     �a@      &@     �D@              Y@      &@      1@      @      @      @      @      @      @                      @      �?              $@             �T@       @      3@      @      @      @      @       @      @                       @              @      .@      �?      *@               @      �?       @                      �?      P@       @      F@       @      (@      �?      @              @      �?      @      �?      @              @@      �?      @@                      �?      4@             �Z@      4@     �J@      @     �B@       @     �@@       @       @              ?@       @      ,@              1@       @      �?              0@       @      @       @      @                       @      *@              @              0@      @               @      0@       @      "@              @       @               @      @             �J@      ,@     �H@      ,@      8@      �?      1@              @      �?              �?      @              9@      *@      @      "@              �?      @       @      @      �?              �?      @               @      @      �?      �?              �?      �?              �?      @              @      �?      @      �?       @              �?      4@      @      (@               @      @      @      @      �?      @      �?       @               @      @              @              @              6@      3@      *@      3@              @      *@      .@      @               @      .@      �?      .@              .@      �?              @              "@             �O@      C@     �F@      C@      F@      C@              @      F@      A@      @      &@       @      &@      �?      @      �?       @               @      �?                      @      �?      @              @      �?              �?             �D@      7@      9@      @      3@       @      "@       @      @       @       @       @              �?       @      �?       @                      �?      �?              @              $@              @      @              �?      @      @      0@      1@      0@      ,@      @      @       @      @              @       @      @              @       @              �?      �?      �?                      �?      *@      @      @              @      @      @      @      @      @      @                      @              @      @                      @      �?              2@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�)�rhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B@D         d                    �?��ے@R�?�           @�@               %                    �?�1�d��?�             l@                                    �?8�Z$���?2            �S@              	                   �-@����>4�?%             L@                                H�%@      �?             @        ������������������������       �                     �?                                83C6@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        
                           �?D>�Q�?"             J@                               ��:3@�>4և��?             <@                                �%@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @                                hލC@���N8�?             5@                                    �?z�G�z�?             @                                 �G@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     0@                                ��|$@r�q��?             8@                                  6@      �?	             0@        ������������������������       �                     @                                pF @�	j*D�?             *@                               �&B@"pc�
�?             &@                               ���@����X�?             @        ������������������������       �                     @        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        !       "                    9@���7�?             6@        ������������������������       �                     $@        #       $                 ���&@�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        &       O                    �?6��L��?e            `b@       '       2                     @��-soi�?M            @\@       (       1                    �?����e��?,            �P@       )       *                    �?�O4R���?"            �J@       ������������������������       �                     A@        +       0                   �<@�}�+r��?             3@        ,       -                     �?r�q��?             @        ������������������������       �                      @        .       /                   �7@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     *@        ������������������������       �        
             *@        3       N                 ���4@z�J��?!            �G@       4       I                 P��%@���Q��?             D@       5       6                    0@X�<ݚ�?             ;@        ������������������������       �                     @        7       <                  sW@      �?             8@        8       9                 ���@      �?              @       ������������������������       �                     @        :       ;                   �7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        =       H                    �?     ��?             0@       >       G                 `�("@������?             .@       ?       F                 `�X!@���Q��?             $@       @       E                 @3�@      �?              @       A       B                 �?�@      �?             @        ������������������������       �                     �?        C       D                   �8@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        J       K                    �?$�q-�?
             *@       ������������������������       �                     $@        L       M                 ���0@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        P       Y                     @      �?             A@        Q       X                     �?     ��?             0@       R       S                    �?�q�q�?             "@        ������������������������       �                     @        T       W                     @      �?             @       U       V                 ���`@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        Z       c                    @�<ݚ�?             2@       [       \                 �̼6@      �?             0@        ������������������������       �                     @        ]       ^                    @$�q-�?	             *@        ������������������������       �                      @        _       `                 ��T?@z�G�z�?             @       ������������������������       �                     @        a       b                 pf�C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        e       �                    �?��Ɛ���?'           p~@       f       �                    �?�=��ny�?�            v@       g       �                    �?$�*7��?�            �u@        h       {                     @r�q��?$             R@        i       j                   �9@���@��?            �B@        ������������������������       �                     &@        k       l                 ���,@�	j*D�?             :@        ������������������������       �                     @        m       x                    �?��<b���?             7@       n       o                   �;@@�0�!��?
             1@        ������������������������       �                     �?        p       w                 p�w@      �?	             0@       q       r                 ���<@��S�ۿ?             .@        ������������������������       �                     @        s       v                    @@      �?              @        t       u                 ��`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        y       z                   @B@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        |       }                    5@(N:!���?            �A@        ������������������������       �                     �?        ~       �                    ?@l��\��?             A@              �                   �<@H%u��?             9@       �       �                   �:@�8��8��?             8@        ������������������������       �                     @        �       �                   @<@ףp=
�?             4@       �       �                 ���@�t����?
             1@        ������������������������       �                     @        �       �                   @@"pc�
�?             &@        ������������������������       ����Q��?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        �       �                     �?<�N��?�            Pq@        �       �                    �?�θ�?            �C@       �       �                 `f�D@��R[s�?            �A@       �       �                 ��$:@�q�q�?             ;@        ������������������������       �                     @        �       �                 03k:@և���X�?             5@        ������������������������       �                      @        �       �                   �<@p�ݯ��?             3@        �       �                   �>@r�q��?             @        ������������������������       �                     @        �       �                   �@@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    R@8�Z$���?	             *@       �       �                   �I@�8��8��?             (@        �       �                 `fF<@z�G�z�?             @        �       �                   @G@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    &@l��\��?�            �m@        ������������������������       �                     �?        �       �                     @\ ���?�            �m@        �       �                 `f�)@ �h�7W�?$            �J@        ������������������������       �                     5@        �       �                    =@     ��?             @@       �       �                    �?r�q��?             2@       �       �                   �*@@�0�!��?             1@       �       �                   �;@���!pc�?             &@       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     ,@        �       �                    �?H� ��w�?s             g@        �       �                  ��@�>����?             ;@        ������������������������       �                     .@        �       �                   @'@r�q��?             (@       �       �                    >@"pc�
�?             &@       �       �                   �<@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?P��-�?d            �c@       �       �                 �T�C@�F����?b            @c@       �       �                   @@@ )�y���?\             b@       �       �                   �>@D���ͫ�?C            @Y@       �       �                   �;@0�>���?=            �V@       �       �                   �:@�U�:��?&            �M@       �       �                   �8@h�����?#             L@       �       �                 �1@����?�?            �F@        �       �                   �4@      �?             0@        ������������������������       �                      @        �       �                  s@      �?              @        ������������������������       �                     @        �       �                   �5@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     =@        �       �                 @33@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     @        ������������������������       �                     @@        �       �                   �?@�z�G��?             $@        ������������������������       �                     �?        �       �                   �@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     F@        �       �                    >@�<ݚ�?             "@       �       �                    ;@���Q��?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �:@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?P�~D&�?N            �`@        �       �                     �?��S���?	             .@       �       �                    C@      �?              @        �       �                   �U@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    7@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @������?E            �]@        �       �                    @���N8�?             5@       ������������������������       �                     0@        ������������������������       �                     @        �       �                     �?�q��/��?:            �X@        �       �                    �?���N8�?             5@       �       �                 03�M@z�G�z�?             .@        �       �                 ��9L@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                   �G@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        �                          0@�C��2(�?,            @S@        �                          �?�GN�z�?             6@       �       �                    +@�d�����?             3@        ������������������������       �                      @        �                       ��l#@@�0�!��?             1@        �       �                    3@�q�q�?             "@        ������������������������       �                     @        �       �                    5@      �?             @        ������������������������       �                     �?                                 �7@���Q��?             @        ������������������������       �                      @                              �&B@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                 �?h㱪��?            �K@                             ��A@`Jj��?             ?@       	                        @@@XB���?             =@        
                         ?@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        
             4@                                 A@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     8@        �t�bh�h*h-K ��h/��R�(KMKK��h]�B       �|@     �o@     �J@     �e@      (@     �P@      &@     �F@       @       @              �?       @      �?       @                      �?      "@     �E@      @      7@      @      @              @      @              �?      4@      �?      @      �?      �?              �?      �?                      @              0@      @      4@      @      (@              @      @      "@       @      "@       @      @              @       @       @              @       @                       @      �?      5@              $@      �?      &@      �?                      &@     �D@     �Z@      8@     @V@      �?     @P@      �?      J@              A@      �?      2@      �?      @               @      �?      @      �?                      @              *@              *@      7@      8@      0@      8@      .@      (@      @              (@      (@      �?      @              @      �?       @               @      �?              &@      @      &@      @      @      @      @       @       @       @      �?              �?       @      �?                       @      @                       @      @                      �?      �?      (@              $@      �?       @               @      �?              @              1@      1@      @      *@      @      @              @      @      @      @      �?              �?      @                       @              @      ,@      @      (@      @              @      (@      �?       @              @      �?      @              �?      �?              �?      �?               @             `y@     @T@     @s@     �F@     0s@      E@      N@      (@      =@       @      &@              2@       @              @      2@      @      ,@      @              �?      ,@       @      ,@      �?      @              @      �?       @      �?              �?       @              @                      �?      @       @               @      @              ?@      @              �?      ?@      @      6@      @      6@       @      @              2@       @      .@       @      @              "@       @      @       @      @              @                      �?      "@             �n@      >@      >@      "@      :@      "@      2@      "@      @              (@      "@               @      (@      @      �?      @              @      �?      �?      �?                      �?      &@       @      &@      �?      @      �?       @      �?       @                      �?       @              @                      �?       @              @              k@      5@              �?      k@      4@      I@      @      5@              =@      @      .@      @      ,@      @       @      @       @                      @      @              �?              ,@             �d@      1@      9@       @      .@              $@       @      "@       @      @       @      @                       @      @              �?             �a@      .@     `a@      .@      a@       @     @W@       @     �U@      @      K@      @      K@       @      F@      �?      .@      �?       @              @      �?      @              @      �?              �?      @              =@              $@      �?              �?      $@                      @      @@              @      @              �?      @       @               @      @              F@               @      @       @      @               @       @      �?              @      @              �?      @              @      �?             �X@      B@      @       @      �?      @      �?       @      �?                       @              @      @      �?              �?      @             �V@      <@      @      0@              0@      @             �U@      (@      0@      @      (@      @      @      @      @                      @       @              @       @      @                       @     �Q@      @      1@      @      ,@      @               @      ,@      @      @      @      @              @      @              �?      @       @       @              �?       @               @      �?               @              @             �J@       @      =@       @      <@      �?       @      �?       @                      �?      4@              �?      �?              �?      �?              8@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJX"4qhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B@G         |                 ��%@�3�n��?�           @�@               '                    �?܈=�Z��?�            �q@               &                    �?�q�q�?/            @Q@                                  �?�#}7��?-            �P@                                03�@������?             ;@        ������������������������       �                      @                                pF @z�G�z�?             9@              	                    �?�LQ�1	�?             7@        ������������������������       �                      @        
                          �2@z�G�z�?             .@        ������������������������       �                      @                                  �5@�θ�?
             *@        ������������������������       �                     �?                                   9@r�q��?	             (@        ������������������������       �                     �?                                ���@"pc�
�?             &@        ������������������������       �                     �?                                ���@ףp=
�?             $@        ������������������������       �                      @                                �&B@      �?              @       ������������������������       �؇���X�?             @        ������������������������       �                     �?        ������������������������       �                      @                                  �4@��(\���?             D@                                �Y�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @               %                   @<@�?�|�?            �B@                                 �:@���7�?             6@        ������������������������       �                     @               $                    �?�}�+r��?             3@               !                 ���@�����H�?             "@        ������������������������       �                     @        "       #                   @@z�G�z�?             @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �        
             .@        ������������������������       �                      @        (       )                     �?0��xX��?�            @k@        ������������������������       �                     @        *       5                   �4@@mW���?�            �j@        +       ,                 �?�@������?            �D@       ������������������������       �                     8@        -       .                 pf� @�t����?
             1@        ������������������������       ��q�q�?             @        /       0                     @@4և���?             ,@        ������������������������       �                     @        1       4                    �?ףp=
�?             $@        2       3                 @�"@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        6       e                 @3�@�R����?t            �e@       7       P                   �;@�q�Q�?C             X@        8       O                    �?���Q��?             >@       9       :                 033@X�<ݚ�?             ;@        ������������������������       �                      @        ;       N                   �:@���Q��?             9@       <       C                    �?      �?             8@        =       >                 ���@����X�?             @        ������������������������       �                     @        ?       @                 �&B@      �?             @        ������������������������       �                     �?        A       B                   �8@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        D       G                 ���@������?             1@        E       F                    7@      �?             @        ������������������������       �                      @        ������������������������       �                      @        H       I                 �?$@8�Z$���?	             *@        ������������������������       �                     @        J       M                 �1@����X�?             @        K       L                   �6@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        Q       ^                 �?�@��IF�E�?-            �P@       R       S                 ��@���#�İ?'            �M@        ������������������������       �                     9@        T       ]                   �@�IєX�?             A@        U       Z                 ��L@"pc�
�?             &@       V       Y                   �>@      �?              @        W       X                 �?$@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        [       \                    D@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     7@        _       d                    �?����X�?             @       `       c                   �A@r�q��?             @       a       b                   �?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     �?        f       o                    �?�s�c���?1            @S@        g       h                     @�q�q�?
             (@        ������������������������       �                     @        i       n                    �?�����H�?             "@       j       k                   �>@؇���X�?             @       ������������������������       �                     @        l       m                 `�("@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        p       w                 ���"@����?'            @P@       q       r                    ?@@��8��?             H@       ������������������������       �                     <@        s       v                   @@@P���Q�?             4@        t       u                 ��i @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             2@        x       {                    $@@�0�!��?
             1@        y       z                   �<@�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        }       �                    �?*�V����?           �z@        ~       �                    �?���PL6�?k            �e@               �                 ��.@�nkK�?#             G@        �       �                    �?�<ݚ�?             "@       �       �                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                    �B@        �       �                   �>@��}� �?H            �_@       �       �                     @�q�q�?)             R@        �       �                    @�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        �       �                     @�0u��A�?"             N@       �       �                    �?l��\��?             A@       ������������������������       �                     6@        �       �                 03�a@      �?             (@       �       �                     �?�����H�?             "@        ������������������������       �                     @        �       �                    �?      �?             @        �       �                   �7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ���i@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 ��1@�θ�?             :@        �       �                   �:@�q�q�?             "@        �       �                    9@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?r�q��?             @        ������������������������       �                     @        �       �                   �;@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        	             1@        �       �                 ��Y.@t�6Z���?            �K@        �       �                    ,@�q�q�?             (@       ������������������������       �                     @        ������������������������       �                     @        �       �                    @Du9iH��?            �E@       ������������������������       �                     D@        ������������������������       �                     @        �       �                    �?�P�����?�            �o@        �       �                    �?ڡR����?            �H@       �       �                   �;@և���X�?            �A@        �       �                    8@�	j*D�?             *@       �       �                    �?�q�q�?             @        ������������������������       �                     @        �       �                    .@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?���!pc�?             6@       �       �                     @�t����?	             1@       �       �                     �?     ��?             0@       �       �                 �;|r@����X�?             ,@       �       �                   �B@r�q��?             (@       �       �                 03SA@����X�?             @       �       �                 �ܵ<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                 ���,@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ��hU@z�G�z�?             @        ������������������������       �                     @        �       �                 @�pX@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   @K@X�Cc�?             ,@       �       �                    �?      �?             (@       �       �                 �̾w@�q�q�?             "@       �       �                    )@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �                            �? 9h�H�?}            `i@        �       �                    �?^|�_��?+            �Q@       �       �                   �>@�\��N��?#            �L@       �       �                   �J@">�֕�?            �A@       �       �                 ��$:@r�q��?             8@        ������������������������       �                      @        �       �                 `f�;@�C��2(�?             6@        ������������������������       �                     ,@        �       �                   @=@      �?              @        ������������������������       �                     �?        �       �                   �<@؇���X�?             @       ������������������������       �                     @        �       �                   @>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 `fF<@���|���?             &@       ������������������������       �                     @        �       �                   @>@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?���!pc�?             6@       �       �                    D@r�q��?             2@        �       �                 03U@�q�q�?             "@       �       �                   �=@      �?              @        �       �                   �7@���Q��?             @        ������������������������       �                     �?        �       �                   �@@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        �       �                 ���[@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �B@����X�?             ,@        �       �                 0�:P@z�G�z�?             @        ������������������������       �                      @        �       �                    �?�q�q�?             @       �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@                                 @fP*L��?R            �`@                                 @�����?             3@       ������������������������       �                     &@                                 @      �?              @       ������������������������       �                     @                                 @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        	                      �T�I@ d�=��?G            @\@       
                        �*@Pa�	�?>            �X@                              ��Y)@�˹�m��?             C@        ������������������������       �                     @                                 @@��a�n`�?             ?@        ������������������������       �                     *@                                �F@r�q��?	             2@                               @D@�q�q�?             "@                               @B@����X�?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                     "@        ������������������������       �        )            �N@                              p�O@X�Cc�?	             ,@                                 ;@      �?              @        ������������������������       �                      @                                 >@      �?             @       ������������������������       ����Q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h*h-K ��h/��R�(KMKK��h]�B�       �{@     �p@     `m@      J@      G@      7@      F@      7@      @      4@       @              @      4@      @      4@               @      @      (@               @      @      $@      �?               @      $@              �?       @      "@      �?              �?      "@               @      �?      @      �?      @              �?       @             �B@      @      �?       @      �?                       @      B@      �?      5@      �?      @              2@      �?       @      �?      @              @      �?      �?      �?      @              $@              .@               @             �g@      =@      @              g@      =@     �C@       @      8@              .@       @       @      �?      *@      �?      @              "@      �?       @      �?       @                      �?      @             @b@      ;@     @S@      3@      2@      (@      .@      (@               @      .@      $@      .@      "@       @      @              @       @       @      �?              �?       @      �?                       @      *@      @       @       @       @                       @      &@       @      @              @       @      �?       @               @      �?              @                      �?      @             �M@      @     �L@       @      9@              @@       @      "@       @      @      �?       @      �?              �?       @              @               @      �?              �?       @              7@               @      @      �?      @      �?       @              �?      �?      �?              @      �?             @Q@       @       @      @              @       @      �?      @      �?      @               @      �?              �?       @               @             �N@      @     �G@      �?      <@              3@      �?      �?      �?              �?      �?              2@              ,@      @      @      @      @                      @       @             `j@     �j@      A@     `a@       @      F@       @      @      �?      @              @      �?              �?       @      �?                       @             �B@      @@     �W@      8@      H@      �?      &@              &@      �?              7@     �B@      @      ?@              6@      @      "@      �?       @              @      �?      @      �?      �?      �?                      �?               @       @      �?       @                      �?      4@      @      @      @       @      �?              �?       @              �?      @              @      �?       @               @      �?              1@               @     �G@      @      @              @      @              @      D@              D@      @              f@     �R@      =@      4@      4@      .@      @      "@      @       @      @              �?       @               @      �?                      @      0@      @      (@      @      &@      @      $@      @      $@       @      @       @      �?       @      �?                       @      @              @                       @      �?      �?              �?      �?              �?              @      �?      @              �?      �?              �?      �?              "@      @      "@      @      @      @      @      �?              �?      @                       @      @                       @     �b@     �K@     �B@      A@      ;@      >@      &@      8@      @      4@       @               @      4@              ,@       @      @      �?              �?      @              @      �?      �?      �?                      �?      @      @      @              �?      @              @      �?              0@      @      .@      @      @      @      @       @      @       @      �?               @       @       @                       @      @                      �?      "@              �?      @      �?                      @      $@      @      �?      @               @      �?       @      �?      �?      �?                      �?              �?      "@             �[@      5@      @      *@              &@      @       @      @              �?       @               @      �?             @Z@       @      X@      @     �A@      @      @              <@      @      *@              .@      @      @      @      @       @      @       @      �?              �?      �?      "@             �N@              "@      @      @      @               @      @      @      @       @              �?      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ;�3whG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM5huh*h-K ��h/��R�(KM5��h|�B@M         �                     @(����7�?�           @�@               !                    �?���}��?�            0t@                                   �?�nkK�?]            @a@                                 �;@0x�!���?P            �]@                                   �?�L���?            �B@                                   �?P���Q�?             4@       ������������������������       �                     *@               	                    )@؇���X�?             @        ������������������������       �                     @        
                          �7@      �?             @        ������������������������       �                      @                                  �8@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   :@�t����?             1@       ������������������������       �        
             ,@                                ��m1@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                  �H@����ȫ�?5            �T@       ������������������������       �        /            �R@                                   �?؇���X�?             @                                   J@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                    �?�KM�]�?             3@                               ���`@؇���X�?             ,@       ������������������������       �        	             &@                                   �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        "       I                    �?p'����?w             g@        #       >                     �?�Gi����?            �B@       $       9                    �?�P�*�?             ?@       %       &                   �3@8����?             7@        ������������������������       �                     �?        '       8                    �?���!pc�?             6@       (       3                  �}S@ҳ�wY;�?             1@       )       *                 �ܵ<@      �?             $@        ������������������������       �                     @        +       2                   �L@����X�?             @       ,       1                    >@r�q��?             @       -       .                   �;@      �?             @        ������������������������       �                     �?        /       0                 03SA@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        4       5                   �?@؇���X�?             @        ������������������������       �                     @        6       7                 �;|r@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        :       ;                   �5@      �?              @        ������������������������       �                     �?        <       =                 @�pX@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ?       H                    �?�q�q�?             @       @       G                    �?z�G�z�?             @       A       B                   �9@      �?             @        ������������������������       �                     �?        C       F                    �?�q�q�?             @       D       E                 ���,@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        J       [                    ,@�V���1�?\            �b@        K       X                   �M@      �?              H@       L       M                     �?����?�?            �F@        ������������������������       �                     @        N       W                    �?�Ń��̧?             E@       O       P                    �?��Y��]�?            �D@        ������������������������       �                     �?        Q       R                 `f�)@�(\����?             D@        ������������������������       �                     .@        S       T                    @@`2U0*��?             9@       ������������������������       �        	             .@        U       V                   @B@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     �?        Y       Z                   �P@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        \       w                   �?@ �o_��?<             Y@       ]       ^                    #@X�Emq�?!            �J@        ������������������������       �                     $@        _       v                    �?�^�����?            �E@       `       m                     �?��i#[�?             E@       a       h                 `fF<@
;&����?             7@       b       g                   �J@�q�q�?
             .@       c       d                   �?@      �?             $@        ������������������������       �                     @        e       f                   �9@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        i       j                   @>@      �?              @        ������������������������       �                      @        k       l                   �J@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        n       o                   �7@�}�+r��?             3@        ������������������������       �                     @        p       q                    �?@4և���?	             ,@       ������������������������       �                     @        r       u                    C@؇���X�?             @        s       t                   �<@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        x       y                    �?�*/�8V�?            �G@        ������������������������       �        
             0@        z       �                    �?�חF�P�?             ?@       {       �                 ���L@��<b���?             7@       |       �                   �C@�q�q�?             (@       }       �                    �?      �?              @        ~                           7@      �?             @        ������������������������       �                     �?        �       �                 `fFJ@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                     �?      �?             @        ������������������������       �                     �?        �       �                    +@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�C��2(�?             &@       ������������������������       �                      @        �       �                �G�:@@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?�e��t�?�            Px@        �       �                    �?@lܯ ��?I            �]@       �       �                    A@�\��N��?-             S@       �       �                   �9@���Q��?)            @P@       �       �                    �?���Q��?            �A@       �       �                    �?��
ц��?             :@        �       �                 ���%@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    -@���Q��?             4@        ������������������������       �                     �?        �       �                    1@p�ݯ��?             3@        ������������������������       �                     @        �       �                    @��S���?             .@        ������������������������       �                      @        �       �                 ���@�n_Y�K�?
             *@        ������������������������       �                     @        �       �                    �?      �?             $@        �       �                   �5@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 �[$@      �?              @       �       �                   �7@և���X�?             @       �       �                    4@�q�q�?             @        �       �                 ��!@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 �̜!@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        �       �                    �?r�q��?             >@        ������������������������       �        
             .@        �       �                   �;@�q�q�?
             .@        �       �                 pf(@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?X�<ݚ�?             "@       �       �                 `�X!@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                   #@�C��2(�?             &@        ������������������������       �                      @        �       �                    I@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?��V#�?            �E@        �       �                    @b�2�tk�?             2@       �       �                 03�-@������?	             .@        �       �                 ��*@      �?              @       �       �                   �;@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �>@H%u��?             9@       �       �                    @���}<S�?             7@       �       �                    �?�t����?             1@       �       �                     @ףp=
�?             $@       �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    #@؇���X�?             @        ������������������������       �                     @        �       �                  `/@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                 `f68@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?PN��T'�?�            �p@        �       �                   @@r֛w���?             ?@        �       �                   @<@      �?	             0@       �       �                    �?�����H�?             "@       �       �                 ���@؇���X�?             @       ������������������������       �                     @        �       �                    9@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?��S���?
             .@       �       �                    �?�n_Y�K�?             *@       �       �                    �?�q�q�?             (@       �       �                   �<@����X�?             @        ������������������������       �                     @        �       �                    ?@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    3@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       4                   @\Qׯ�?�            �m@       �       �                    @%4 �?�            `l@        �       �                    �?z�G�z�?             $@        �       �                 03�;@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       3                0�H@T���.�?�             k@       �       �                   �2@�S	���?�            `j@        ������������������������       �                     ?@        �       2                ���!@ףp=
�?v            �f@       �       1                   �?d/�@7�?]             a@       �       0                @Q!@     ��?X             `@              /                  @F@�? Da�?W            �_@                                �?Ԫ2��?P            �\@                                �:@�����H�?             2@        ������������������������       �                     @                                �=@؇���X�?
             ,@                             03�@z�G�z�?             $@        ������������������������       �                      @        ������������������������       �      �?              @        ������������������������       �                     @        	                      �?�@8��8���?C             X@       
                      �1@@4և���?*             L@                                =@(N:!���?            �A@                                7@�<ݚ�?             2@                                �5@ףp=
�?             $@                                �4@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @                                �8@      �?              @        ������������������������       �                     �?                                �:@����X�?             @        ������������������������       �                      @                              �?$@���Q��?             @                             03s@�q�q�?             @        ������������������������       �                     �?                              ��@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     1@        ������������������������       �                     5@              &                @3�@      �?             D@               %                  �D@     ��?             0@       !      "                  �:@X�Cc�?             ,@        ������������������������       �                     @        #      $                  �A@�eP*L��?             &@       ������������������������       �      �?             @        ������������������������       ����Q��?             @        ������������������������       �                      @        '      .                ��y @      �?             8@       (      )                   4@�S����?             3@        ������������������������       ��q�q�?             @        *      -                   =@      �?             0@       +      ,                ��) @$�q-�?
             *@       ������������������������       �        	             (@        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     (@        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                    �E@        ������������������������       �                     @        ������������������������       �                     (@        �t�b�      h�h*h-K ��h/��R�(KM5KK��h]�BP       �{@      q@      b@     @f@      @     �`@      @     �\@      @      A@      �?      3@              *@      �?      @              @      �?      @               @      �?      �?      �?                      �?       @      .@              ,@       @      �?              �?       @              �?     @T@             �R@      �?      @      �?       @      �?                       @              @       @      1@       @      (@              &@       @      �?              �?       @                      @     `a@      G@      6@      .@      2@      *@      0@      @              �?      0@      @      &@      @      @      @      @               @      @      �?      @      �?      @              �?      �?       @               @      �?                       @      �?              @      �?      @               @      �?       @                      �?      @               @      @      �?              �?      @              @      �?              @       @      @      �?      @      �?      �?               @      �?      �?      �?              �?      �?              �?              �?                      �?     @]@      ?@     �F@      @      F@      �?      @             �D@      �?      D@      �?      �?             �C@      �?      .@              8@      �?      .@              "@      �?              �?      "@              �?              �?       @               @      �?              R@      <@      >@      7@              $@      >@      *@      =@      *@      &@      (@      $@      @      @      @      @               @      @       @                      @      @              �?      @               @      �?      @              @      �?              2@      �?      @              *@      �?      @              @      �?       @      �?       @                      �?      @              �?              E@      @      0@              :@      @      2@      @       @      @      @      @       @       @      �?              �?       @      �?                       @       @       @              �?       @      �?              �?       @              @              $@      �?       @               @      �?              �?       @               @             pr@     �W@     @P@      K@      B@      D@      :@     �C@      5@      ,@      (@      ,@      @       @               @      @               @      (@      �?              @      (@              @      @       @       @              @       @              @      @      @      �?      �?      �?                      �?      @      @      @      @       @      @      �?       @      �?                       @      �?       @               @      �?              �?              �?              "@              @      9@              .@      @      $@      �?      @              @      �?              @      @      @      @      @                      @               @      $@      �?       @               @      �?       @                      �?      =@      ,@      @      &@      @      &@      @      @      �?      @              @      �?              @                      @      @              6@      @      5@       @      .@       @      "@      �?      @      �?              �?      @               @              @      �?      @               @      �?              �?       @              @              �?      �?              �?      �?             �l@      D@      7@       @      .@      �?       @      �?      @      �?      @              �?      �?      �?                      �?       @              @               @      @       @      @      @      @      @       @      @               @       @               @       @               @      @              @       @              �?                       @     �i@      @@     `h@      @@       @       @       @      @              @       @                      @      h@      8@      h@      2@      ?@             @d@      2@     �]@      2@     �[@      2@     �[@      0@     �X@      0@      0@       @      @              (@       @       @       @       @              @       @      @             �T@      ,@      J@      @      ?@      @      ,@      @      "@      �?      @      �?      @                      �?      @              @      @              �?      @       @       @              @       @      �?       @              �?      �?      �?      �?                      �?       @              1@              5@              >@      $@      "@      @      "@      @      @              @      @      @      @      @       @               @      5@      @      0@      @      �?       @      .@      �?      (@      �?      (@                      �?      @              @              (@                       @      "@             �E@                      @      (@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�3hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B@G         |                     @(����7�?�           @�@                                   /@�Ҹf���?�             t@        ������������������������       �                     8@                                   �?P�]���?�            �r@                                   �?�94�s0�?H            �\@                                  �?��v$���?&            �N@                                 �G@��Y��]�?            �D@       ������������������������       �                    �A@        	       
                 ���;@r�q��?             @        ������������������������       �                     @                                ,w�U@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     4@                                   �?�X�<ݺ?"             K@                                 �;@Du9iH��?            �E@                                    �?z�G�z�?	             .@                                   �?���Q��?             @        ������������������������       �                      @                                   5@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                   �?ףp=
�?             $@        ������������������������       �                     @                                  �9@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     <@        ������������������������       �                     &@               {                 @�:x@�s�;�w�?t            �f@              \                     �?DG��L�?r            �f@                7                    �?��+7��?8             W@        !       0                    �?8^s]e�?             =@       "       /                 ���S@8����?             7@       #       .                    �?��S���?	             .@       $       -                 @�6M@�n_Y�K�?             *@       %       ,                    A@���!pc�?             &@       &       +                    ?@և���X�?             @       '       *                    =@z�G�z�?             @       (       )                 �ܵ<@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        1       6                    �?�q�q�?             @       2       3                    �?z�G�z�?             @        ������������������������       �                      @        4       5                    6@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        8       [                    �?���N8�?&            �O@       9       Z                    R@���3�E�?              J@       :       Y                 03�U@ \� ���?            �H@       ;       T                    �?��[�p�?            �G@       <       M                   �>@�I�w�"�?             C@       =       >                 ��I/@�q�q�?             8@        ������������������������       �                     @        ?       L                   �L@X�<ݚ�?             2@       @       E                    @@և���X�?	             ,@        A       D                   �<@      �?             @       B       C                 `fF<@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        F       G                 03k:@�z�G��?             $@        ������������������������       �                      @        H       K                   `H@      �?              @       I       J                   �F@և���X�?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        N       S                   @B@@4և���?             ,@       O       P                   �A@      �?              @        ������������������������       �                     @        Q       R                 ��yC@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        U       V                   @K@�����H�?             "@        ������������������������       �                     @        W       X                 `f�N@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     &@        ]       f                   �?@����!p�?:             V@       ^       e                    &@���J��?#            �I@        _       `                    @@4և���?             ,@        ������������������������       �                     @        a       d                   �6@ףp=
�?             $@        b       c                   �1@      �?             @        ������������������������       �                      @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                    �B@        g       v                    �?������?            �B@       h       u                    �? 	��p�?             =@       i       l                   @A@@4և���?             <@        j       k                 `fF)@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        m       t                   �*@`2U0*��?             9@       n       s                   �F@�IєX�?	             1@        o       p                   �'@؇���X�?             @        ������������������������       �                      @        q       r                   @D@z�G�z�?             @        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     $@        ������������������������       �                      @        ������������������������       �                     �?        w       z                   �:@      �?              @        x       y                   �@@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        }       �                    �?R�}e�.�?�            `x@        ~       �                    �?X�'����?G             _@              �                  ��@և���X�?9            �X@        �       �                 03�@x�����?            �C@        ������������������������       �                     @        �       �                 ���@4?,R��?             B@        ������������������������       �        	             3@        �       �                 0�w@�t����?             1@       �       �                    �?�q�q�?             .@       �       �                   �5@�z�G��?             $@        ������������������������       �                      @        �       �                    9@      �?              @        ������������������������       �                     @        ������������������������       �z�G�z�?             @        �       �                    4@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�Ƀ aA�?#            �M@        �       �                  S�-@�\��N��?             3@        �       �                 Ь* @ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     "@        �       �                 P��%@      �?             D@        �       �                    �?�S����?             3@       �       �                   �8@z�G�z�?	             .@        ������������������������       �                     "@        �       �                 @3�@      �?             @        ������������������������       �                     �?        �       �                   �>@���Q��?             @        ������������������������       �                      @        �       �                  SE"@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 03�1@և���X�?             5@       �       �                   �D@d}h���?             ,@       �       �                    �?8�Z$���?             *@        ������������������������       �                     @        �       �                     @z�G�z�?             $@       �       �                    +@����X�?             @        ������������������������       �                     @        �       �                   �0@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �@@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    @ȵHPS!�?             :@       �       �                    @�IєX�?
             1@        ������������������������       �                     �?        ������������������������       �        	             0@        �       �                    @�<ݚ�?             "@        ������������������������       �                     @        �       �                    @���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �                       �T�I@�{�@�N�?�            �p@       �       �                    �?>a�����?�            �o@        �       �                   @@\X��t�?             7@       �       �                    9@z�G�z�?	             $@        �       �                 ��y@�q�q�?             @        ������������������������       �                     �?        �       �                 ���@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ���@؇���X�?             @        ������������������������       �                      @        �       �                   @<@z�G�z�?             @       ������������������������       �      �?             @        ������������������������       �                     �?        �       �                 83##@�n_Y�K�?             *@        �       �                    @@      �?             @       �       �                   �<@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?����X�?             @       �       �                 `v�0@�q�q�?             @        ������������������������       �                     �?        �       �                   �2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �                          @X�
����?�             m@       �       �                 @3�@�r�.kx�?�            @j@       �       �                 �?�@�{��?��?E             [@       �       �                   �;@�C��2(�?=             V@        �       �                    �?�MI8d�?            �B@       �       �                   �:@r�q��?             >@       �       �                   �4@ �Cc}�?             <@        ������������������������       �        	             ,@        �       �                 ��L@d}h���?
             ,@       �       �                   �8@�q�q�?             "@        �       �                 ���@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?؇���X�?             @       �       �                 ��@z�G�z�?             @        ������������������������       �                     @        �       �                 �&B@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?`'�J�?#            �I@        �       �                  s�@r�q��?	             (@        ������������������������       �                     @        �       �                    >@      �?              @        �       �                   �<@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �C@        �       �                    �?�z�G��?             4@       �       �                   �A@@�0�!��?             1@       �       �                    �?�z�G��?             $@       �       �                   �:@և���X�?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �                          �?�v�\�?>            �Y@       �                         �0@��.N"Ҭ?*            @Q@        �                        �̌!@r�q��?             @       ������������������������       �z�G�z�?             @        ������������������������       �                     �?                                �<@ ������?'            �O@       ������������������������       �                    �D@                                 �?���7�?             6@                             ���"@�X�<ݺ?             2@       ������������������������       �                     1@        ������������������������       �                     �?        ������������������������       �                     @        	                      ��Y7@6YE�t�?            �@@       
                         �?���N8�?             5@                                 �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?                                 %@������?             .@        ������������������������       �                     @        ������������������������       �        	             &@        ������������������������       �                     (@                                 @���7�?             6@                              ���A@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             0@                                 @�eP*L��?             &@                                ;@�q�q�?             "@        ������������������������       �                      @                                 >@և���X�?             @       ������������������������       ����Q��?             @        ������������������������       �                      @        ������������������������       �                      @        �t�bh�h*h-K ��h/��R�(KMKK��h]�B�       �{@      q@     `c@     �d@              8@     `c@     �a@      @     �[@      �?      N@      �?      D@             �A@      �?      @              @      �?      �?      �?                      �?              4@      @     �I@      @      D@      @      (@       @      @               @       @      �?              �?       @              �?      "@              @      �?      @              @      �?                      <@              &@     �b@      @@     �b@      =@      Q@      8@      4@      "@      0@      @       @      @       @      @       @      @      @      @      @      �?      @      �?      @                      �?      �?                       @      @                       @               @       @              @       @      @      �?       @               @      �?              �?       @                      �?      H@      .@     �B@      .@     �B@      (@     �B@      $@      =@      "@      0@       @      @              $@       @      @       @      @      �?       @      �?       @                      �?      �?              @      @               @      @      @      @      @       @      @      �?                      �?      @              *@      �?      @      �?      @               @      �?              �?       @              @               @      �?      @              @      �?              �?      @                       @              @      &@             �T@      @      I@      �?      *@      �?      @              "@      �?      @      �?       @              �?      �?      @             �B@             �@@      @      ;@       @      :@       @       @      �?      �?              �?      �?      8@      �?      0@      �?      @      �?       @              @      �?      @              �?      �?      $@               @              �?              @       @      �?       @               @      �?              @                      @     �q@     @Z@     @P@     �M@      E@      L@       @      ?@      @              @      ?@              3@      @      (@      @      $@      @      @       @              �?      @              @      �?      @       @      @       @                      @               @      A@      9@      "@      $@      "@      �?              �?      "@                      "@      9@      .@      0@      @      (@      @      "@              @      @              �?      @       @       @              �?       @               @      �?              @              "@      (@      @      &@       @      &@              @       @       @       @      @              @       @       @       @                       @              @      �?              @      �?      @                      �?      7@      @      0@      �?              �?      0@              @       @      @              @       @               @      @             �k@      G@     �j@      D@      *@      $@       @       @       @      �?      �?              �?      �?              �?      �?              @      �?       @              @      �?      @      �?      �?              @       @      @      @      �?      @      �?                      @       @               @      @       @      �?      �?              �?      �?      �?                      �?              @     @i@      >@     �f@      =@     �U@      6@      T@       @      ?@      @      9@      @      9@      @      ,@              &@      @      @      @      �?      @      �?                      @      @              @                       @      @      �?      @      �?      @              �?      �?              �?      �?               @             �H@       @      $@       @      @              @       @       @       @       @      �?              �?      @             �C@              @      ,@      @      ,@      @      @      @      @      �?               @      @              @              @      @             �W@      @     �P@       @      @      �?      @      �?      �?              O@      �?     �D@              5@      �?      1@      �?      1@                      �?      @              <@      @      0@      @      @      �?      @                      �?      &@      @              @      &@              (@              5@      �?      @      �?              �?      @              0@              @      @      @      @               @      @      @      @       @               @       @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ� �NhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B�F         j                    �?�6��l�?�           @�@               i                    @f����?�            �p@              ^                   �>@>���Rp�?�            Pp@              !                     @�7�?r            �g@                                03�a@�8��8��?1             U@                                   �?hA� �?)            �Q@        ������������������������       �                     =@                                   6@��p\�?            �D@       	                          �1@��2(&�?             6@       
                           �?�X�<ݺ?             2@                                  �?�IєX�?             1@                               ��Y)@      �?
             0@        ������������������������       �                     @                                   �?ףp=
�?             $@        ������������������������       �                      @                                   :@      �?              @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?                                    @      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     3@                                   �?����X�?             ,@        ������������������������       �                     @                                   �?և���X�?             @        ������������������������       �                     �?                                   �8@�q�q�?             @                                   @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        "       ;                    �?�G��l��?A            @Z@        #       :                    @p9W��S�?             C@       $       -                    �?V������?            �B@        %       (                 03�-@��S���?	             .@       &       '                 P��+@�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        )       ,                 ���.@r�q��?             @        *       +                   �<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        .       9                    �?"pc�
�?             6@       /       0                   �0@؇���X�?
             5@        ������������������������       �                     @        1       8                    �?r�q��?	             2@       2       3                    7@      �?             (@        ������������������������       �                     �?        4       7                 `f�@"pc�
�?             &@       5       6                  s�@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       ������H�?             "@        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        <       ]                 ��Y1@�#}7��?,            �P@       =       T                 `f�%@z�J��?            �G@       >       S                    ;@      �?             @@       ?       @                    $@��
ц��?             :@        ������������������������       �                     @        A       B                 ���@�eP*L��?             6@        ������������������������       �                     @        C       R                    �?X�<ݚ�?             2@       D       Q                   �9@      �?
             0@       E       P                    �?����X�?	             ,@       F       O                    7@�q�q�?             (@       G       N                 �[$@      �?              @       H       K                    4@և���X�?             @        I       J                 ��!@      �?             @        ������������������������       �                      @        ������������������������       �                      @        L       M                 �̜!@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        U       V                    �?������?	             .@       ������������������������       �                      @        W       X                    +@և���X�?             @        ������������������������       �                      @        Y       \                    �?z�G�z�?             @       Z       [                    ;@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     4@        _       h                    �?�k~X��?1             R@        `       g                    �?P���Q�?             4@       a       f                    �?�X�<ݺ?
             2@        b       e                 ��T@؇���X�?             @        c       d                   �G@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                      @        ������������������������       �        &             J@        ������������������������       �                      @        k       t                    *@2�Bo��?(           �{@        l       m                     @)O���?             B@        ������������������������       �                     &@        n       s                     @`�Q��?             9@        o       p                   X1@�����H�?             "@       ������������������������       �                     @        q       r                 pf�3@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     0@        u       �                    �?B�a���?           py@       v       �                    �?ɍo�?�            �t@       w       �                 ��$:@h~��M�?�            �t@       x       �                 ���+@����x9�?�            �p@       y       �                 ��\+@(��Le�?�            �m@       z                           �?l��\��?�            �m@        {       |                   �<@ �q�q�?             8@       ������������������������       �                     2@        }       ~                   �=@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?��hq��?�            �j@        �       �                    >@ȵHPS!�?             :@       �       �                   �<@@�0�!��?             1@       �       �                  s�@��S�ۿ?             .@        ������������������������       �                     @        �       �                 ��(@�����H�?             "@       ������������������������       �؇���X�?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     "@        �       �                 ���$@�B!A�?{            �g@       �       �                   �>@�Km�a̾?]            �a@       �       �                     @(;L]n�?=            �V@        ������������������������       �                     @        �       �                 ��@XB���?:            �U@        ������������������������       �                      @        �       �                   �:@`��>�ϗ?8            @U@       ������������������������       �                    �I@        �       �                 pb@г�wY;�?             A@        �       �                 ��@r�q��?             @       ������������������������       �                     @        �       �                   �;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     <@        �       �                 �&B@H%u��?              I@        ������������������������       �                     0@        �       �                   �@@�0�!��?             A@        �       �                    D@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 �?�@��� ��?             ?@        ������������������������       �                     "@        �       �                   �?@"pc�
�?             6@        ������������������������       �                     �?        �       �                   �B@؇���X�?             5@       �       �                 @3�@$�q-�?             *@        ������������������������       �                     @        �       �                 pF� @ףp=
�?             $@       �       �                   �@@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                 @3�@      �?              @        ������������������������       ��q�q�?             @        ������������������������       �                     @        �       �                    &@r�q��?             H@        �       �                   @H@�θ�?             *@       �       �                   �5@ףp=
�?	             $@        �       �                   �1@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                     @        �       �                   �P@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �;@؇���X�?            �A@        ������������������������       �                     *@        �       �                 `f�)@�GN�z�?             6@        ������������������������       �                     @        �       �                    =@�d�����?             3@        �       �                   �*@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    @@�r����?	             .@        ������������������������       �                     @        �       �                   �F@"pc�
�?             &@       �       �                   @D@����X�?             @       �       �                   @B@r�q��?             @       ������������������������       �      �?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     >@        �       �                   �F@Ɣ��Hr�?#            �M@       �       �                    ?@      �?             C@       �       �                   `@@8����?             7@        �       �                   �<@��
ц��?             *@       �       �                 �ܵ<@�z�G��?             $@       �       �                 ��";@���Q��?             @       ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@        �       �                 0��F@z�G�z�?	             .@       �       �                    <@      �?              @        ������������������������       �                     @        �       �                    �?���Q��?             @       �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?��s����?             5@       �       �                    �?�<ݚ�?
             2@        �       �                 �̬L@؇���X�?             @       �       �                   �L@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                 �T@@���!pc�?             &@       �       �                    R@      �?              @       �       �                    K@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �                           �?�=A�F�?=             S@        �       �                    �?� �	��?             9@        �       �                 p"�X@      �?              @       �       �                    �?r�q��?             @       �       �                   �:@z�G�z�?             @        ������������������������       �                     @        �       �                 ��hU@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    9@ҳ�wY;�?             1@        ������������������������       �                     @        �                         �C@և���X�?             ,@        �                           �?z�G�z�?             @       �       �                   @K@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @                              ���[@�<ݚ�?             "@       ������������������������       �                     @                                  @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                �:@�:�]��?)            �I@                                ?@������?            �B@       	                        �9@@4և���?             <@        
                      ���@z�G�z�?             $@        ������������������������       �                     @                                 �?����X�?             @        ������������������������       �                     �?                                 �?r�q��?             @                              hfF#@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     2@                                 �?�<ݚ�?             "@                                 @�q�q�?             @                                 C@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     ,@        �t�bh�h*h-K ��h/��R�(KMKK��h]�B�       0{@     Pq@     �Q@     �h@     �O@     �h@      O@     �_@      @     @S@      @     �P@              =@      @      C@      @      3@      �?      1@      �?      0@      �?      .@              @      �?      "@               @      �?      @      �?       @              @              �?              �?       @       @       @                       @              3@      @      $@              @      @      @              �?      @       @      �?       @      �?                       @      @             �K@      I@      &@      ;@      &@      :@      @       @      @      @              @      @              �?      @      �?       @      �?                       @              @      @      2@      @      2@              @      @      .@      @      "@      �?               @      "@      �?      "@              �?      �?       @      �?                      @      �?                      �?      F@      7@      8@      7@      4@      (@      ,@      (@      @              $@      (@              @      $@       @      $@      @      $@      @       @      @      @      @      @      @       @       @       @                       @      �?       @               @      �?              �?              @               @                       @               @      @              @      &@               @      @      @               @      @      �?      @      �?      @                      �?      �?              4@              �?     �Q@      �?      3@      �?      1@      �?      @      �?       @               @      �?                      @              &@               @              J@       @             �v@     �S@      1@      3@              &@      1@       @      �?       @              @      �?       @      �?                       @      0@             �u@      N@     �q@     �F@     �q@     �F@     �n@      6@      k@      6@      k@      5@      7@      �?      2@              @      �?              �?      @             @h@      4@      7@      @      ,@      @      ,@      �?      @               @      �?      @      �?       @                       @      "@             `e@      1@     ``@      "@     �U@      @      @              U@      @               @      U@      �?     �I@             �@@      �?      @      �?      @              �?      �?              �?      �?              <@              F@      @      0@              <@      @      �?       @               @      �?              ;@      @      "@              2@      @              �?      2@      @      (@      �?      @              "@      �?       @      �?              �?       @              �?              @       @      �?       @      @              D@       @      $@      @      "@      �?       @      �?      �?              �?      �?      @              �?       @               @      �?              >@      @      *@              1@      @      @              ,@      @      �?      @              @      �?              *@       @      @              "@       @      @       @      @      �?      @      �?       @                      �?      @                      �?      >@              B@      7@      3@      3@      0@      @      @      @      @      @      @       @      �?       @       @                      @      @              $@              @      (@      @      @              @      @       @       @       @               @       @              �?                      @      1@      @      ,@      @      @      �?       @      �?              �?       @              @               @      @      @      @      @      �?              �?      @                       @      @              @              @             �N@      .@      ,@      &@      @      @      �?      @      �?      @              @      �?      �?      �?                      �?              �?       @              &@      @      @               @      @      �?      @      �?       @      �?                       @               @      @       @      @              �?       @               @      �?             �G@      @     �@@      @      :@       @       @       @      @              @       @              �?      @      �?       @      �?              �?       @              @              2@              @       @      @       @      �?       @               @      �?              @              @              ,@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ���bhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM7huh*h-K ��h/��R�(KM7��h|�B�M         x                     @\H�l�?�           @�@               M                     �?,siC��?�            �r@              L                    @�G�z��?g             d@              9                    �?H���I�?f            �c@                                  �?�ϡz�?D            �[@                                03[=@���N8�?             E@                                  �H@�q�q�?             @        ������������������������       �                     @        	       
                    K@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     B@               8                   �L@<��¤�?)             Q@              '                   �@@     8�?&             P@              &                 0�/[@">�֕�?            �A@              %                    �?��>4և�?             <@                               �ܵ<@��}*_��?             ;@                                �̌*@"pc�
�?             &@        ������������������������       �                     @                                   �?����X�?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @                                   �?      �?             0@                                03SA@�q�q�?             @        ������������������������       �                     @                                  �;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @               $                   �<@���Q��?             $@              #                 `f�D@և���X�?             @                                  `@@z�G�z�?             @        ������������������������       �                      @        !       "                   �A@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        (       )                   @B@П[;U��?             =@        ������������������������       �                     @        *       +                   @E@\X��t�?             7@        ������������������������       �                     @        ,       -                    �?j���� �?
             1@        ������������������������       �                      @        .       7                    �?��S���?	             .@       /       6                 `f�;@և���X�?             ,@       0       5                   �J@z�G�z�?             $@       1       4                   �G@�����H�?             "@        2       3                 ��:@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        :       ;                    �?r�qG�?"             H@       ������������������������       �                     9@        <       G                 Ј�V@\X��t�?             7@       =       @                    �?      �?             0@        >       ?                 ��+T@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        A       F                    D@"pc�
�?
             &@        B       E                    �?      �?             @       C       D                   �B@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        H       I                   �E@؇���X�?             @        ������������������������       �                     @        J       K                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        N       ]                   �'@nIz~]�?\            �a@        O       \                    &@����>�?            �B@       P       Y                   @E@�4�����?             ?@       Q       R                    �?z�G�z�?             9@        ������������������������       �                     @        S       T                    @�C��2(�?             6@        ������������������������       �                     @        U       X                   �6@�����H�?             2@        V       W                   �1@����X�?             @        ������������������������       �                      @        ������������������������       ����Q��?             @        ������������������������       �                     &@        Z       [                   �P@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ^       _                    .@��
P��?H            @Z@        ������������������������       �        	             (@        `       a                    �?�P�*�??            @W@        ������������������������       �                    �A@        b       o                 ���+@ 	��p�?&             M@        c       n                 ��\+@H%u��?             9@       d       m                   �*@�8��8��?             8@       e       j                   @D@�C��2(�?             6@       f       i                    =@�X�<ݺ?             2@       g       h                   �;@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@        k       l                   �F@      �?             @        ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        p       q                    �?Pa�	�?            �@@        ������������������������       �        	             ,@        r       s                   �?@�}�+r��?             3@        ������������������������       �                     &@        t       w                   �@@      �?              @        u       v                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        y       .                   @xN�%�F�?           �y@       z       �                    �?V�e��n�?�            Pw@        {       |                    @�b��[��?"            �K@        ������������������������       �                     @        }       �                    �? �o_��?              I@        ~       �                    7@      �?
             ,@               �                    �?      �?             @       �       �                 H�%@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                  S�2@���Q��?             $@       �       �                 H�%@և���X�?             @        ������������������������       �                      @        �       �                    �?z�G�z�?             @       �       �                   �<@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   �7@tk~X��?             B@        �       �                 ��y@և���X�?             @        ������������������������       �                     �?        �       �                    �?�q�q�?             @       �       �                    /@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ��&@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   @<@ܷ��?��?             =@       �       �                   @@؇���X�?             5@       �       �                   �:@d}h���?             ,@        ������������������������       �                     �?        �       �                 ���@�θ�?             *@        ������������������������       �                     @        ������������������������       ��z�G��?             $@        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?��{��2�?�            �s@        �       �                    �?�Q����?0             T@       �       �                    B@^��>�b�?'            @P@       �       �                    �?��Q:��?"            �M@        �       �                 @�@և���X�?	             ,@       �       �                    �?���Q��?             $@       �       �                 ���@      �?              @       �       �                  s�@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �=@�L�lRT�?            �F@       �       �                    @�xGZ���?            �A@       �       �                    �?�ʻ����?             A@       �       �                 P��@��}*_��?             ;@        ������������������������       �                     @        �       �                   �9@�eP*L��?             6@        �       �                 ���/@���!pc�?             &@       �       �                  � @      �?              @       �       �                    4@z�G�z�?             @        ������������������������       �                      @        �       �                   �7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                 `f7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 �?�@"pc�
�?             &@        �       �                    ;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�����H�?             "@       �       �                 @3�@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 pf�3@����X�?             @       �       �                    &@���Q��?             @        ������������������������       �                     �?        �       �                 ���)@      �?             @        ������������������������       �                     �?        �       �                    ;@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     @        �       �                    @�q�q�?	             .@        �       �                   �8@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                 pfv2@�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?��w\ud�?�            �m@        �       �                    �?XB���?             =@       �       �                   �<@ �q�q�?             8@       ������������������������       �                     4@        �       �                   �>@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    &@4�d����?�             j@        ������������������������       �                     @        �       -                �T�E@�d2 Λ�?�            �i@       �                         �<@�
F%u�?�             i@       �                          �?�	a�$a�?U            ``@       �       �                 �1@\����?P            @^@        �       �                    �?b�h�d.�?            �A@       �       �                    4@      �?             @@        ������������������������       �                      @        �       �                 ��@r�q��?             8@        ������������������������       �                     �?        �       �                 ���@�LQ�1	�?             7@       �       �                 ���@��S�ۿ?             .@        �       �                    7@r�q��?             @        ������������������������       �                     @        �       �                   �8@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        �       �                   �5@      �?              @        ������������������������       �                     �?        �       �                    :@؇���X�?             @        ������������������������       �                     @        �       �                 �?$@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        �       �                   �7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �                         �4@��+��<�?7            �U@                               ��Y @�C��2(�?             6@                              �?�@z�G�z�?             $@        ������������������������       �                     @                                 �?����X�?             @                               �1@r�q��?             @        ������������������������       �                      @        ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                     (@        	      
                pf� @     ��?)             P@       ������������������������       �                    �E@                                 �?���N8�?             5@                               �;@@4և���?             ,@                                �9@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     @        ������������������������       �                     $@              "                  @@@�~t��?.            @Q@                                �=@���|���?             6@                              ���"@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                �>@�����?	             3@        ������������������������       �                     @                                �?@���Q��?             .@                              pff@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @                                �@      �?              @        ������������������������       �                     �?               !                @3�@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        #      $                �?�@`�q�0ܴ?#            �G@        ������������������������       �                     7@        %      ,                   �?�8��8��?             8@       &      +                   �?�KM�]�?             3@       '      *                @3�@؇���X�?             ,@        (      )                  �D@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �        
             &@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        /      6                   @@-�_ .�?            �B@        0      1                   @�<ݚ�?             "@       ������������������������       �                     @        2      3                   @�q�q�?             @        ������������������������       �                     �?        4      5                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     <@        �t�b��     h�h*h-K ��h/��R�(KM7KK��h]�Bp       �|@     �o@     `a@     `d@      M@     �Y@      L@     �Y@     �E@     �P@       @      D@       @      @              @       @      �?       @                      �?              B@     �D@      ;@     �B@      ;@      8@      &@      1@      &@      1@      $@      "@       @      @              @       @      �?              @       @       @       @       @      @              @       @      �?              �?       @              @      @      @      @      �?      @               @      �?       @      �?                       @       @              @                      �?      @              *@      0@              @      *@      $@      @              @      $@               @      @       @      @       @       @       @      �?       @      �?       @      �?                       @              @      �?              @              �?              @              *@     �A@              9@      *@      $@      (@      @      @       @               @      @              "@       @       @       @       @      �?       @                      �?              �?      @              �?      @              @      �?      �?      �?                      �?       @             @T@     �N@      ;@      $@      5@      $@      4@      @              @      4@       @      @              0@       @      @       @       @              @       @      &@              �?      @              @      �?              @              K@     �I@              (@      K@     �C@             �A@      K@      @      6@      @      6@       @      4@       @      1@      �?       @      �?       @                      �?      "@              @      �?      �?      �?       @               @                      �?      @@      �?      ,@              2@      �?      &@              @      �?      �?      �?              �?      �?              @             �s@      W@     �q@     �V@      B@      3@              @      B@      ,@      @      @      @      �?       @      �?              �?       @              �?              @      @      @      @               @      @      �?       @      �?       @                      �?       @                      @      =@      @      @      @      �?               @      @      �?      @      �?                      @      �?      �?      �?                      �?      :@      @      2@      @      &@      @      �?              $@      @      @              @      @      @               @             �n@     �Q@      C@      E@      <@     �B@      6@     �B@      @       @      @      @      @      @      �?      @      �?                      @      @               @                      @      0@      =@      0@      3@      .@      3@      $@      1@              @      $@      (@       @      @      @      �?      @      �?       @               @      �?              �?       @              @              �?       @               @      �?               @      "@      �?      �?              �?      �?              �?       @      �?      @              @      �?                      @      @       @      @       @              �?      @      �?      �?               @      �?       @                      �?       @              �?                      $@      @              $@      @      @       @      @                       @      @      @              @      @              j@      =@      <@      �?      7@      �?      4@              @      �?              �?      @              @             �f@      <@              @     �f@      7@     �f@      3@     �^@      "@      \@      "@      =@      @      <@      @       @              4@      @              �?      4@      @      ,@      �?      @      �?      @               @      �?              �?       @              "@              @       @              �?      @      �?      @              @      �?       @      �?      �?              �?       @      �?                       @     �T@      @      4@       @       @       @      @              @       @      @      �?       @              @      �?              �?      (@             �O@      �?     �E@              4@      �?      *@      �?      @      �?      @                      �?      $@              @              $@             �M@      $@      ,@       @      �?       @      �?                       @      *@      @      @              "@      @      @      @      @                      @      @       @              �?      @      �?      @                      �?     �F@       @      7@              6@       @      1@       @      (@       @      �?       @      �?      �?              �?      &@              @              @                      @     �A@       @      @       @      @              �?       @              �?      �?      �?      �?                      �?      <@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ+�MhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM)huh*h-K ��h/��R�(KM)��h|�B@J         B                    �?�JX-��?�           @�@               1                    �?      �?O            �^@                                  �?4��@���??             Y@                                   �?��P���?            �D@              
                   �G@�q�q�?             8@                                   @�}�+r��?             3@       ������������������������       �                     .@               	                 ���%@      �?             @       ������������������������       �                     @        ������������������������       �                     �?                                ,w�U@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?                                    @������?             1@       ������������������������       �                     *@        ������������������������       �                     @               $                     �?0B��D�?'            �M@                                  �:@�G�z��?             4@                                  �5@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @                                ��hU@����X�?	             ,@                                  @@"pc�
�?             &@                                  �?�<ݚ�?             "@                               03SA@����X�?             @                               �ܵ<@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @                !                    �?�q�q�?             @        ������������������������       �                     �?        "       #                   �H@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        %       ,                   �7@8�Z$���?            �C@        &       '                 ��y@      �?              @        ������������������������       �                     �?        (       )                    5@����X�?             @        ������������������������       �                     @        *       +                 ���@      �?             @        ������������������������       �                      @        ������������������������       �                      @        -       .                 83�0@�g�y��?             ?@       ������������������������       �                     :@        /       0                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        2       3                 03�-@���|���?             6@        ������������������������       �                     @        4       9                    �?@�0�!��?             1@       5       6                 ��U@�C��2(�?             &@       ������������������������       �                     @        7       8                    F@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        :       A                 Ј�_@�q�q�?             @       ;       <                     @z�G�z�?             @        ������������������������       �                      @        =       @                    @�q�q�?             @       >       ?                   �<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        C       �                    �?J,K/c�?w           p�@        D       Q                     @4��PH��?y            �g@       E       F                    �?�*v��?=            @X@       ������������������������       �                     G@        G       P                   �;@�t����?            �I@        H       K                   �8@      �?             8@       I       J                 ���`@�X�<ݺ?	             2@       ������������������������       �                     1@        ������������������������       �                     �?        L       M                    �?r�q��?             @        ������������������������       �                     @        N       O                     �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     ;@        R       c                   �5@�\@k!�?<            �V@        S       V                 03�@r�q��?             8@        T       U                 ��}@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        W       \                    �?��2(&�?             6@        X       Y                    �?�q�q�?             @        ������������������������       �                      @        Z       [                    @      �?             @        ������������������������       �                      @        ������������������������       �                      @        ]       b                    @      �?
             0@        ^       _                    @r�q��?             @        ������������������������       �                     @        `       a                 ��T?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        d       �                 @3�2@�2�,��?,            �P@       e       p                    �?*;L]n�?&             N@        f       g                    9@�z�G��?             4@        ������������������������       �                     @        h       o                    �?ҳ�wY;�?             1@       i       n                    �?     ��?
             0@       j       k                 ���@X�Cc�?             ,@        ������������������������       �                     @        l       m                 `f�@"pc�
�?             &@       ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        q       �                 P��%@      �?             D@       r       s                    @`�Q��?             9@        ������������������������       �                     @        t       �                    �?�GN�z�?             6@       u       �                    K@���N8�?             5@       v       �                 `��!@z�G�z�?             4@       w       �                 `�X!@      �?             0@       x                          �;@z�G�z�?             .@       y       ~                   �9@      �?             @       z       }                 pff@      �?             @        {       |                   �7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?z�G�z�?             .@       �       �                    �?���!pc�?             &@       �       �                    D@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �/@��v����?�             y@       �       �                   @N@���T��?�            �o@       �       �                    �?Xa9g�U�?�             o@       �       �                     @@Ix�<��?�            �m@        �       �                    @XB���?              M@        ������������������������       �                     *@        �       �                   �*@`Ӹ����?            �F@       �       �                   �<@P���Q�?             D@       �       �                   �(@�8��8��?             8@       �       �                    &@��S�ۿ?             .@       �       �                   �5@�8��8��?             (@        �       �                   �1@r�q��?             @        ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �:@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        
             0@        ������������������������       �                     @        �       �                 ��@�3�۸��?z            `f@        �       �                 ���@����X�?             @       �       �                    �?r�q��?             @        ������������������������       �                     �?        �       �                 ���	@z�G�z�?             @       �       �                   �B@      �?             @       �       �                    6@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 �?�@���@�c�?t            �e@       �       �                    �? r���??            �W@        �       �                   �=@���N8�?             5@       �       �                  ��@�IєX�?             1@        ������������������������       �                     @        �       �                 ��(@ףp=
�?             $@       ������������������������       ������H�?             "@        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �?@`׀�:M�?2            �R@       ������������������������       �        &             L@        �       �                   @@@�X�<ݺ?             2@        �       �                   �@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        
             0@        �       �                   @@@�C��2(�?5            @S@       �       �                    �?�����H�?(             K@        ������������������������       �                     �?        �       �                   �<@���C��?'            �J@       �       �                   �0@@4և���?             E@        �       �                 pFD!@z�G�z�?             @        ������������������������       �      �?              @        ������������������������       �                     @        �       �                   �9@@-�_ .�?            �B@        ������������������������       �                     0@        �       �                   �;@�����?             5@        ������������������������       �                     �?        �       �                 ��) @P���Q�?             4@        ������������������������       �                     &@        �       �                 pf� @�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �>@���!pc�?	             &@        �       �                   �=@z�G�z�?             @        �       �                 �̌!@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �?@�q�q�?             @        ������������������������       �                     �?        �       �                 ��I @z�G�z�?             @       ������������������������       �      �?             @        ������������������������       �                     �?        �       �                   �E@�nkK�?             7@       ������������������������       �        	             0@        �       �                   �F@؇���X�?             @        �       �                 @3�@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        �       �                 hfF"@      �?             @        ������������������������       �                     �?        �       �                   �P@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       (                  �R@�Ҳ���?Y            �b@       �       !                   �?`K�����?X            @b@       �                           @�t����?H            �]@       �                          �?�Sb(�	�?@             [@       �                         �J@V�a�� �?#             M@       �       �                 ��$:@������?            �F@        ������������������������       �                     (@        �       �                   �>@���|���?            �@@        �       �                   �E@�z�G��?             $@        ������������������������       �                     @        �       �                   �=@���Q��?             @       �       �                   �F@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     �?        �                          �?��<b���?             7@       �       �                     @���N8�?             5@       �       �                 ��yC@@4և���?             ,@        �       �                 �TaA@z�G�z�?             @        ������������������������       �                     @        �       �                   @B@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        �                           >@և���X�?             @       ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     *@                                 �?z�):���?             I@                             ���0@�eP*L��?             F@        ������������������������       �                     @                                 ,@�n_Y�K�?            �C@        ������������������������       �                     @        	                         D@���!pc�?            �@@       
                          �?$��m��?             :@                                 <@؇���X�?             @        ������������������������       �                     @                                �@@      �?             @        ������������������������       �                     �?        ������������������������       �                     @                                  @�S����?	             3@                               �7@�θ�?             *@        ������������������������       �                     @                                �?@      �?              @        ������������������������       �                     @                                �@@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                                 L@      �?             @                                )@      �?             @        ������������������������       �                      @                                 :@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     &@        "      '                pf�C@ 7���B�?             ;@        #      $                ��T?@�C��2(�?             &@       ������������������������       �                     "@        %      &                   @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             0@        ������������������������       �                     @        �t�bh�h*h-K ��h/��R�(KM)KK��h]�B�       @}@     �n@     �N@     �N@     �J@     �G@      "@      @@      @      3@      �?      2@              .@      �?      @              @      �?              @      �?      @                      �?      @      *@              *@      @              F@      .@      &@      "@      �?      @      �?                      @      $@      @      "@       @      @       @      @       @       @       @       @                       @      @               @               @              �?       @              �?      �?      �?              �?      �?             �@@      @      @      @      �?               @      @              @       @       @               @       @              >@      �?      :@              @      �?              �?      @               @      ,@      @              @      ,@      �?      $@              @      �?      @              @      �?               @      @      �?      @               @      �?       @      �?      �?      �?                      �?              �?      �?             py@     �f@     �M@      `@      @     �V@              G@      @     �F@      @      2@      �?      1@              1@      �?              @      �?      @               @      �?       @                      �?              ;@     �J@      C@      4@      @      �?      �?      �?                      �?      3@      @      @       @       @               @       @               @       @              .@      �?      @      �?      @              �?      �?      �?                      �?      $@             �@@      A@      :@      A@      @      ,@              @      @      &@      @      &@      @      "@      @               @      "@              "@       @                       @      �?              4@      4@      1@       @              @      1@      @      0@      @      0@      @      (@      @      (@      @      @      @      @      �?      �?      �?              �?      �?               @                       @      "@                      �?      @                      �?      �?              @      (@      @       @      �?       @               @      �?               @                      @      @             �u@      K@     �m@      .@     �m@      *@      l@      *@      L@       @      *@             �E@       @      C@       @      6@       @      ,@      �?      &@      �?      @      �?      @               @      �?      @              @               @      �?       @                      �?      0@              @              e@      &@      @       @      @      �?      �?              @      �?      @      �?      �?      �?      �?                      �?       @              �?                      �?     `d@      "@     @W@       @      4@      �?      0@      �?      @              "@      �?       @      �?      �?              @             @R@      �?      L@              1@      �?      �?      �?              �?      �?              0@             �Q@      @      H@      @      �?             �G@      @     �C@      @      @      �?      �?      �?      @             �A@       @      0@              3@       @              �?      3@      �?      &@               @      �?              �?       @               @      @      @      �?       @      �?       @                      �?       @              @       @              �?      @      �?      @      �?      �?              6@      �?      0@              @      �?      �?      �?              �?      �?              @              (@               @       @      �?              �?       @               @      �?             �[@     �C@     �[@      B@      U@     �A@     @R@     �A@      G@      (@     �@@      (@      (@              5@      (@      @      @              @      @       @      @      �?       @      �?      �?                      �?      2@      @      0@      @      *@      �?      @      �?      @              �?      �?              �?      �?              "@              @      @      @      �?              @       @              *@              ;@      7@      8@      4@              @      8@      .@              @      8@      "@      1@      "@      �?      @              @      �?      @      �?                      @      0@      @      $@      @      @              @      @      @              �?      @              @      �?              @              @              @      @      �?      @               @      �?      �?      �?                      �?       @              &@              :@      �?      $@      �?      "@              �?      �?              �?      �?              0@                      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJY]hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM=huh*h-K ��h/��R�(KM=��h|�B@O         T                    �?��!h
��?�           @�@               G                 p�H@>��C��?�             m@                                   @l��
I��?m            @d@                                   6@hA� �?+            �Q@                                  �?�L���?            �B@                                 �2@�#-���?            �A@                               `f�)@�IєX�?             A@        ������������������������       �                     ,@        	                          �*@ףp=
�?             4@       
                           :@�r����?             .@        ������������������������       ����Q��?             @        ������������������������       �                     $@        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                    �@@               &                    �?I� ��?B             W@                                03�@����>�?            �B@        ������������������������       �                      @               %                 ��.@4�2%ޑ�?            �A@                                  1@l��
I��?             ;@        ������������������������       �                     @               "                    �?�ՙ/�?             5@                                 �5@�θ�?	             *@        ������������������������       �                     �?                                   �?r�q��?             (@        ������������������������       �                     �?                                   9@"pc�
�?             &@        ������������������������       �                     �?                                 ��@z�G�z�?             $@        ������������������������       �                     �?                !                 ���@�����H�?             "@        ������������������������       �                     �?        ������������������������       �      �?              @        #       $                   �<@      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        '       0                   �3@���|���?*            �K@        (       )                 �"-@X�<ݚ�?             2@        ������������������������       �                      @        *       +                    �?z�G�z�?	             $@        ������������������������       �                     �?        ,       -                 ��T?@�<ݚ�?             "@       ������������������������       �                     @        .       /                    @      �?             @        ������������������������       �                      @        ������������������������       �                      @        1       F                    �?����>�?            �B@       2       A                 ���.@J�8���?             =@       3       @                    �?�q�q�?             8@       4       9                   �9@j���� �?             1@        5       8                 pff@�����H�?             "@        6       7                   �7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        :       ;                 ��Y@      �?              @        ������������������������       �                     �?        <       =                   �;@؇���X�?             @        ������������������������       �                     @        >       ?                 ��� @      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        B       C                    ;@���Q��?             @        ������������������������       �                     �?        D       E                     @      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        H       I                    �?��?^�k�?+            �Q@       ������������������������       �        #            �L@        J       S                    @8�Z$���?             *@       K       R                    �?�8��8��?             (@       L       M                    �?�����H�?             "@        ������������������������       �                      @        N       Q                   @B@؇���X�?             @       O       P                 ���`@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        U       �                     �?�q�q�?5            ~@        V       ]                   �;@T��o��?A            @W@        W       X                    �?�z�G��?             $@        ������������������������       �                     @        Y       Z                    �?      �?             @        ������������������������       �                      @        [       \                 �̰f@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ^       {                    �?̠�4��?9            �T@        _       z                   �M@� �	��?             9@       `       s                   �H@�û��|�?             7@       a       b                 ���<@X�<ݚ�?             2@        ������������������������       �                     @        c       f                 `f�A@��S���?             .@        d       e                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        g       h                   �?@���Q��?             $@        ������������������������       �                      @        i       j                   �A@      �?              @        ������������������������       �                     �?        k       n                    �?և���X�?             @        l       m                 @�Cq@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        o       p                   @H@�q�q�?             @        ������������������������       �                     �?        q       r                 ���X@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        t       y                    �?z�G�z�?             @       u       x                 �D8H@      �?             @       v       w                 ��L@@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        |       �                    @>���Rp�?&             M@       }       �                   �J@^(��I�?%            �K@       ~       �                    >@�X����?             F@               �                 `fF:@�S����?             3@        ������������������������       �                     @        �       �                 `fF<@�θ�?	             *@        ������������������������       �                     �?        �       �                 `f�D@r�q��?             (@       �       �                   �A@      �?              @       �       �                   �<@؇���X�?             @       �       �                   �>@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?� �	��?             9@       �       �                    �?�û��|�?             7@       �       �                 ��I/@���|���?             6@        ������������������������       �                     @        �       �                 03k:@D�n�3�?             3@        ������������������������       �                     @        �       �                    �?     ��?             0@       �       �                   �G@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        �       �                    �?      �?             @       �       �                 03�Q@      �?             @        ������������������������       �                      @        �       �                   �D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �                     @        �       �                    �?T������?�            0x@        �       �                 ���@@��x_F-�?!            �I@       �       �                 ؼC1@r�q��?             H@       �       �                     @z�G�z�?             D@        �       �                 `��,@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 033.@��G���?            �B@       �       �                    +@r�q��?             B@        ������������������������       �                      @        �       �                    ?@�t����?             A@       �       �                   �<@r�q��?             8@       �       �                    �?�LQ�1	�?             7@       �       �                   @@�S����?             3@       �       �                 ��y@z�G�z�?             .@        ������������������������       �                     �?        �       �                 ���@d}h���?             ,@        �       �                    9@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    5@z�G�z�?             $@        ������������������������       �                     �?        �       �                    9@�����H�?             "@        ������������������������       �                     @        �       �                   @<@r�q��?             @       ������������������������       �z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                      @        �       �                    *@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    !@i#[�G�?�             u@        �       �                     @�û��|�?             7@        ������������������������       �                      @        �       �                    @���Q��?
             .@       �       �                 ���8@��
ц��?	             *@        ������������������������       �                     @        �       �                    �?�z�G��?             $@       ������������������������       �                     @        �       �                 ��T?@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                     @@�y����?�            �s@        �       �                    �?�IєX�?+             Q@       �       �                   @F@ ,��-�?&            �M@       �       �                    �?dP-���?            �G@       �       �                   �3@������?            �D@       �       �                    C@      �?             @@       �       �                    @��a�n`�?             ?@        ������������������������       �                     @        �       �                 `fF)@H%u��?             9@        �       �                    &@ףp=
�?             $@       �       �                   �5@      �?              @        �       �                   �1@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   �;@�r����?	             .@       ������������������������       �                     &@        �       �                    ?@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     @        ������������������������       �        	             (@        ������������������������       �                     "@        �       8                �T�I@ZՏ�m|�?�            �n@       �                         �;@�+����?�            `m@        �                       �1@H�V�e��?=            �Y@        �       �                    �?�99lMt�?            �C@        ������������������������       �                      @        �       �                 �?$@؀�:M�?            �B@       �       �                    �?�θ�?             :@       �       �                    7@���N8�?             5@       ������������������������       �        	             ,@        �       �                   �8@����X�?             @        ������������������������       �                      @        �       �                   �:@���Q��?             @       �       �                 ���@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �7@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �5@���!pc�?             &@        ������������������������       �                     @                                 �9@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @                                �:@�����H�?&            �O@                                �?85�}C�?%            �N@                             ��Y @ i���t�?            �H@                                �?�חF�P�?             ?@             
                  �3@\-��p�?             =@              	                �?�@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     7@                                 �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     2@        ������������������������       �                     (@        ������������������������       �                      @              3                   �?ՀJ��?W            �`@                                �?HVĮ���?S            �_@                                 �?�����?             5@                               �<@�t����?             1@       ������������������������       �                     "@                                 >@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @              2                   �?�NW���?F            �Z@                             �?�@<����?>            �W@       ������������������������       �        !             G@              1                   �?ZՏ�m|�?            �H@             $                @3�@�㙢�c�?             G@               !                  �?@      �?             $@        ������������������������       �                      @        "      #                  �A@      �?              @        ������������������������       �                     @        ������������������������       ����Q��?             @        %      0                  �=@�8��8��?             B@       &      -                  �<@��2(&�?             6@       '      ,                  @<@�IєX�?
             1@       (      +                pf� @��S�ۿ?	             .@        )      *                ��) @z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                      @        .      /                ���"@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        	             ,@        ������������������������       �                     @        ������������������������       �                     &@        4      5                �ܭ2@�q�q�?             @        ������������������������       �                     @        6      7                   �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        9      <                p�O@�z�G��?             $@       :      ;                   >@      �?              @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                      @        �t�bh�h*h-K ��h/��R�(KM=KK��h]�B�       �z@     �q@      I@     �f@      H@     �\@      @     �P@      @      A@      @      @@       @      @@              ,@       @      2@       @      *@       @      @              $@              @      �?                       @             �@@     �F@     �G@      $@      ;@       @               @      ;@       @      3@              @       @      *@      @      $@      �?               @      $@              �?       @      "@              �?       @       @      �?              �?       @              �?      �?      @      @      @      @                      @               @     �A@      4@       @      $@               @       @       @      �?              @       @      @               @       @               @       @              ;@      $@      3@      $@      1@      @      $@      @       @      �?      �?      �?              �?      �?              @               @      @      �?              �?      @              @      �?      @      �?                      @      @               @      @      �?              �?      @              @      �?               @               @      Q@             �L@       @      &@      �?      &@      �?       @               @      �?      @      �?       @               @      �?                      @              @      �?             �w@      Y@     �N@      @@      @      @              @      @      @       @              �?      @              @      �?              M@      9@      ,@      &@      ,@      "@      $@       @      @              @       @      �?      @              @      �?              @      @       @              @      @              �?      @      @      @      �?      @                      �?      �?       @              �?      �?      �?              �?      �?              @      �?      @      �?      �?      �?      �?                      �?       @              �?                       @      F@      ,@     �D@      ,@      >@      ,@      0@      @      @              $@      @              �?      $@       @      @       @      @      �?      @      �?              �?      @               @                      �?      @              ,@      &@      ,@      "@      ,@       @      @              &@       @              @      &@      @       @       @       @                       @      @      @      �?      @               @      �?      �?              �?      �?               @                      �?               @      &@              @             �s@      Q@     �D@      $@      D@       @      @@       @       @      �?              �?       @              >@      @      >@      @               @      >@      @      4@      @      4@      @      0@      @      (@      @      �?              &@      @      @      �?              �?      @               @       @              �?       @      �?      @              @      �?      @      �?      �?              @              @                      �?      $@                      �?       @              �?       @               @      �?             `q@      M@      "@      ,@               @      "@      @      @      @              @      @      @      @              �?      @      �?                      @       @             �p@      F@      P@      @     �K@      @     �E@      @     �B@      @      <@      @      <@      @      @              6@      @      "@      �?      @      �?       @      �?       @                      �?      @               @              *@       @      &@               @       @              �?       @      �?              �?      "@              @              (@              "@             �i@      D@     @i@     �@@     @T@      5@      9@      ,@       @              7@      ,@      4@      @      0@      @      ,@               @      @               @       @      @       @       @               @       @                      �?      @      �?      @                      �?      @       @              @      @      @      @                      @      L@      @      L@      @      F@      @      :@      @      9@      @       @      @       @                      @      7@              �?      �?              �?      �?              2@              (@                       @     @^@      (@     @]@      $@      3@       @      .@       @      "@              @       @               @      @              @             �X@       @     �U@       @      G@             �D@       @      C@       @      @      @               @      @      @      @               @      @     �@@      @      3@      @      0@      �?      ,@      �?      @      �?      @                      �?      $@               @              @       @      @                       @      ,@              @              &@              @       @      @              �?       @               @      �?              @      @      �?      @      �?      �?              @       @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ4
hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B�G         T                    �?������?�           @�@               	                     @��1+�?�            �m@                                  �H@�Ru߬Α?L            �\@       ������������������������       �        B            @Y@                                   �?$�q-�?
             *@                                   J@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        
       ?                    �?l��TO��?L            @_@              >                   �A@�L�lRT�?5            �V@              =                 03�7@��i#[�?2             U@                               03�@d�� z�?0            @T@        ������������������������       �                      @               <                    @ܩ�d	��?/            �S@              '                    �?��Sݭg�?.            �S@               &                    �?r�q��?             E@              !                    �?>A�F<�?             C@                                 �0@     ��?             @@        ������������������������       �                     @                                   �?�+e�X�?             9@                                  �6@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                  �5@��<b���?             7@        ������������������������       �                     �?                                   9@"pc�
�?
             6@        ������������������������       �                     �?                                ���@��s����?	             5@        ������������������������       �                      @                                 pF @�KM�]�?             3@       ������������������������       �                     1@        ������������������������       �                      @        "       %                    �?r�q��?             @        #       $                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        (       )                 �&B@*O���?             B@        ������������������������       �                     "@        *       ;                 P��%@|��?���?             ;@       +       :                    �?�����?             3@       ,       3                 @3�@ҳ�wY;�?             1@        -       2                 �?�@և���X�?             @       .       /                    4@      �?             @        ������������������������       �                      @        0       1                    ;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        4       9                   �>@z�G�z�?             $@       5       8                    3@�����H�?             "@        6       7                  �M$@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        @       M                    �?4�2%ޑ�?            �A@        A       B                 ��"@��
ц��?
             *@        ������������������������       �                     @        C       H                   �;@�z�G��?	             $@       D       G                    @؇���X�?             @       E       F                 `f7@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        I       J                  S�2@�q�q�?             @        ������������������������       �                     �?        K       L                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        N       O                 ��T?@���7�?             6@       ������������������������       �                     ,@        P       S                    @      �?              @       Q       R                 ��p@@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        U       X                    @�Sn��?*           �}@        V       W                    @�q�q�?	             .@       ������������������������       �                     $@        ������������������������       �                     @        Y       �                 ��i=@�n�vb&�?!           �|@       Z       �                    �?t��I��?�            Pv@       [       �                   �F@�e��[�?�            �r@       \       w                    �? �L�T�?�            @o@        ]       ^                 ���@�'�`d�?            �@@        ������������������������       �                     @        _       f                     @R�}e�.�?             :@        `       a                   �9@      �?              @        ������������������������       �                     @        b       e                    =@z�G�z�?             @       c       d                 ���,@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        g       n                   @@�q�q�?             2@       h       i                    5@�<ݚ�?             "@        ������������������������       �                     �?        j       k                    9@      �?              @        ������������������������       �                      @        l       m                   @<@r�q��?             @       ������������������������       �z�G�z�?             @        ������������������������       �                     �?        o       t                   �<@X�<ݚ�?             "@       p       q                 `v�0@z�G�z�?             @        ������������������������       �                     @        r       s                   �2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        u       v                    @@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        x       �                 ��$:@TW@k��?�             k@       y       �                    �?\�sl���?�            �j@       z       �                 �{@�`�k�?�             j@        {       �                    �?r�q��?9            �V@        |       }                  s�@�8��8��?             8@        ������������������������       �                      @        ~       �                    >@      �?             0@              �                   �<@r�q��?             (@       �       �                 ��(@�C��2(�?             &@       ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                     @F.< ?�?)            �P@        ������������������������       �                     "@        �       �                 ���@�MWl��?#            �L@       �       �                 ��@��� ��?             ?@        �       �                 ��@      �?              @       �       �                  ��	@z�G�z�?             @       �       �                   �>@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    B@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 ���@�nkK�?             7@        �       �                 ���@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     .@        �       �                 �?$@$��m��?             :@        �       �                   �7@���Q��?             $@        ������������������������       �                     @        �       �                   �=@և���X�?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        �       �                    >@     ��?             0@       �       �                   �8@8�Z$���?             *@       �       �                 �1@ףp=
�?             $@        �       �                   �5@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   �;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                 `fF)@T(y2��?K            �]@       �       �                   �B@ p�/��?:            @V@       �       �                 ���!@��Y��]�?5            �T@       �       �                 @Q!@�&=�w��?$            �J@       �       �                   �>@p���?!             I@       ������������������������       �                     B@        �       �                   �?@@4և���?	             ,@        ������������������������       �                     �?        ������������������������       �                     *@        �       �                    8@�q�q�?             @        ������������������������       �                     �?        �       �                   �;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     =@        �       �                 @3�@����X�?             @       �       �                   �D@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                     @�r����?             >@       �       �                    @@PN��T'�?             ;@       ������������������������       �                     1@        �       �                   @A@���Q��?             $@        ������������������������       �                     @        �       �                   �3@؇���X�?             @       �       �                   @D@z�G�z�?             @        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                 03k:@���Q��?             @        ������������������������       �                     �?        �       �                   @B@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     G@        �       �                    5@��GEI_�?"            �N@        �       �                    �?�θ�?             *@        �       �                   �2@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                    @      �?              @        �       �                 �!4@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?@��8��?             H@       �       �                    �?������?             B@       ������������������������       �                     >@        �       �                    :@r�q��?             @        ������������������������       �                     @        �       �                 ��,/@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     (@        �                       �̾w@@VK��\�?B            @Y@       �                          �?�Y �K�?@            @X@       �                        D�_@hP�vCu�?6            �T@       �                        D�\@��J�fj�?1            �R@       �                           �?���Q��?0            �Q@       �       �                   �D@T�7�s��?&            �L@       �       �                    �?��
ц��?            �C@       �       �                 `f�A@�\��N��?             3@        �       �                    �?z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        �       �                 0w�W@�<ݚ�?             "@       �       �                    �?      �?              @        �       �                   �;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   @B@�G�z��?
             4@       �       �                   �;@X�Cc�?             ,@        �       �                 8�T@      �?              @       �       �                    6@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       	                   �?�<ݚ�?             2@       �                         �J@�z�G��?             $@       �       �                    �?؇���X�?             @        ������������������������       �                      @                                 �H@z�G�z�?             @                             ���X@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                 �?�q�q�?             @                             ��L@@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        
                        �H@      �?              @        ������������������������       �                     @                                 @@      �?             @                                �J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @                                 �?�θ�?
             *@        ������������������������       �                     @                                pA@�z�G��?             $@        ������������������������       �                     @                                 �?և���X�?             @                                >@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?                                 +@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        
             .@        ������������������������       �                     @        �t�b�      h�h*h-K ��h/��R�(KMKK��h]�B�        |@     `p@      N@     `f@      �?     @\@             @Y@      �?      (@      �?      @      �?                      @              "@     �M@     �P@      @@      M@      :@      M@      7@      M@       @              5@      M@      4@      M@      @     �A@      @      ?@      @      :@              @      @      3@      �?      �?      �?                      �?      @      2@      �?              @      2@              �?      @      1@       @               @      1@              1@       @              �?      @      �?      �?      �?                      �?              @              @      *@      7@              "@      *@      ,@      *@      @      &@      @      @      @      @      �?       @              �?      �?              �?      �?                      @       @       @       @      �?      �?      �?              �?      �?              @                      �?       @                       @      �?              @              @              ;@       @      @      @      @              @      @      �?      @      �?      @              @      �?                      �?       @      �?      �?              �?      �?              �?      �?              5@      �?      ,@              @      �?      @      �?              �?      @              �?             `x@     �T@      @      $@              $@      @             x@     @R@      t@     �B@     pp@     �@@      k@     �@@      :@      @      @              3@      @      @      �?      @              @      �?      @      �?              �?      @              �?              (@      @      @       @              �?      @      �?       @              @      �?      @      �?      �?              @      @      @      �?      @              �?      �?      �?                      �?      �?      @              @      �?             �g@      :@     �g@      7@     @g@      7@     �R@      .@      6@       @       @              ,@       @      $@       @      $@      �?      @      �?      @                      �?      @             �J@      *@      "@              F@      *@      ;@      @      @      @      @      �?      @      �?              �?      @              �?              �?       @               @      �?              6@      �?      @      �?      @                      �?      .@              1@      "@      @      @      @              @      @       @      @      �?              &@      @      &@       @      "@      �?       @      �?              �?       @              @               @      �?              �?       @                      @     �[@       @     @U@      @      T@       @     �I@       @     �H@      �?      B@              *@      �?              �?      *@               @      �?      �?              �?      �?              �?      �?              =@              @       @      �?       @      �?      �?              �?      @              :@      @      7@      @      1@              @      @              @      @      �?      @      �?      @              �?      �?       @              @              @               @      @              �?       @       @              �?       @      �?      G@             �L@      @      $@      @      @       @      @                       @      @      �?       @      �?              �?       @              @             �G@      �?     �A@      �?      >@              @      �?      @               @      �?       @                      �?      (@             @P@      B@     @P@      @@      I@      @@      E@      @@      E@      <@      @@      9@      2@      5@      "@      $@       @       @               @       @              @       @      @      �?       @      �?              �?       @              @                      �?      "@      &@      "@      @      @      @      �?      @      �?                      @       @              @                      @      ,@      @      @      @      @      �?       @              @      �?      �?      �?              �?      �?              @              �?       @      �?      �?      �?                      �?              �?      @      �?      @              @      �?      �?      �?              �?      �?               @              $@      @      @              @      @      @              @      @       @      �?       @                      �?       @       @               @       @                      @       @              .@                      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ��;hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B�G         �                 0�&H@\H�l�?�           @�@                                  #@�#�����?d           P�@               
                 03�;@N{�T6�?&            �K@               	                    @ 	��p�?             =@                               P��%@h�����?             <@                                �(\�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     :@        ������������������������       �                     �?                                   @R�}e�.�?             :@                                   !@      �?              @       ������������������������       �                     @        ������������������������       �                      @                                   �?�X�<ݺ?             2@        ������������������������       �                     $@                                ��T?@      �?              @       ������������������������       �                     @                                pf�C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                ���@l���?>           ��@                                    @`���i��?             F@        ������������������������       �                     &@                                P��@Pa�	�?            �@@        ������������������������       �                     0@                                   :@�IєX�?             1@        ������������������������       �                     $@                                   A@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @                [                    �?�Q�9�?(           p~@        !       ,                     @�3[�s(�?`            �b@        "       +                   �;@�1�`jg�?(            �K@        #       *                   �7@R���Q�?             4@        $       %                    �?���!pc�?             &@       ������������������������       �                     @        &       '                    �?      �?             @        ������������������������       �                     �?        (       )                    �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                    �A@        -       Z                 ��Y7@�q���?8             X@       .       W                   �=@\�Uo��?/             S@       /       0                   �-@� ���?)            @P@        ������������������������       �                      @        1       8                 ��@և���X�?'            �O@        2       7                   �5@�KM�]�?
             3@        3       6                    �?����X�?             @        4       5                 03�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     (@        9       V                    @~�4_�g�?             F@       :       E                    �?      �?             D@        ;       D                   �<@X�Cc�?             ,@       <       C                    �?�q�q�?
             (@       =       B                    �?���|���?	             &@       >       A                  S�-@���Q��?             $@        ?       @                 Ь* @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        F       I                   �9@�θ�?             :@        G       H                    �?�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        J       U                    @�q�q�?
             .@       K       R                    �?X�Cc�?	             ,@       L       O                    ;@�q�q�?             "@        M       N                 xF�'@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        P       Q                    �?����X�?             @        ������������������������       �                     @        ������������������������       �                      @        S       T                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        X       Y                   @B@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �        	             4@        \       y                    �?��?"m�?�             u@        ]       x                    �?�q�q��?             H@       ^       u                  I>@�5��
J�?             G@       _       j                 @Q,@RB)��.�?            �E@       `       a                     @8����?             7@        ������������������������       �                      @        b       c                   �7@���N8�?             5@        ������������������������       �                      @        d       i                    =@�S����?             3@       e       f                 ���@      �?             (@       ������������������������       �                     @        g       h                   @@և���X�?             @       ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     @        k       t                    �?ףp=
�?             4@       l       m                   �8@r�q��?             (@        ������������������������       �                     @        n       s                 �ܵ<@�q�q�?             @       o       r                  A7@z�G�z�?             @        p       q                     @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        v       w                 `f�A@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        z       {                 ���@8��8���?�             r@        ������������������������       �                     �?        |       �                     �?4B��@�?�            �q@        }       �                   �Q@�c�Α�?             =@       ~       �                   �>@      �?             <@              �                 `fF<@�q�q�?	             2@       �       �                   �E@�θ�?             *@        ������������������������       �                     �?        �       �                   �G@r�q��?             (@        ������������������������       �                     @        �       �                    J@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �J@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                 �TaA@ףp=
�?             $@        ������������������������       �                     @        �       �                 ��yC@      �?             @        �       �                   @B@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?����"$�?�             p@       �       �                   @N@x�kE�?v            `g@       �       �                     @HKS�l�?s            �f@        �       �                    �?�7��?            �C@        ������������������������       �                      @        �       �                   �*@@-�_ .�?            �B@       �       �                    =@�>����?             ;@        �       �                   �;@؇���X�?             ,@       ������������������������       �                     $@        �       �                   �'@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        	             *@        ������������������������       �                     $@        �       �                 �?�@���Hx�?Z             b@        �       �                   �@P�2E��?)            @P@       �       �                    �?@4և���?             E@        �       �                   �=@@4և���?
             ,@       �       �                  s�@�C��2(�?             &@        ������������������������       �                     @        �       �                 ��(@      �?              @       ������������������������       �؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ���@@4և���?             <@        ������������������������       �                     &@        �       �                    ;@�t����?	             1@       ������������������������       �                     &@        �       �                   �=@�q�q�?             @        ������������������������       �                     �?        �       �                   �?@z�G�z�?             @        ������������������������       �                      @        �       �                    D@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     7@        �       �                    �?p#�����?1            �S@       �       �                    �?$�Z����?/             S@        ������������������������       �                     �?        �       �                 ���!@���?.            �R@       �       �                   �0@����>4�?!             L@        ������������������������       �                     @        �       �                   �2@f1r��g�?             �J@        ������������������������       �                     "@        �       �                   �3@"pc�
�?             F@        ������������������������       ����Q��?             @        �       �                 pf� @8�Z$���?            �C@       �       �                   �>@     ��?             @@       ������������������������       �                     3@        �       �                   �?@�θ�?
             *@        ������������������������       �                     �?        �       �                   �@@r�q��?	             (@        �       �                 @3�@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                 @3�@�����H�?             "@        ������������������������       ��q�q�?             @        ������������������������       �                     @        �       �                    8@և���X�?             @        ������������������������       �                     @        �       �                   �;@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     3@        ������������������������       �                     @        �       �                     @      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                     @0z�(>��?#            �Q@        ������������������������       �        	             .@        �       �                    6@�h����?             L@        �       �                    @�θ�?             *@       �       �                    �?և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                    �E@        �                          @X�Cc�?Q            �_@       �                         �H@$� _��?L            �]@       �                          �?      �?@             Y@       �       �                   �;@��|�5��?<            �W@        �       �                    �?��a�n`�?             ?@        ������������������������       �                     0@        �       �                    �?z�G�z�?
             .@       �       �                    �?ףp=
�?             $@        ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                      @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 `f�K@���Q��?             @        ������������������������       �                     �?        �       �                     @      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �                       03?U@0�� ��?*            �O@       �       �                    �?h+�v:�?             A@        �       �                 `f�L@��
ц��?	             *@       �       �                      @����X�?             @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �z�G�z�?             @        �       �                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�q�q�?             5@       ������������������������       �        	             (@        �                       ЈrS@�<ݚ�?             "@                                @K@      �?             @        ������������������������       �                     �?                                 >@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                 G@V�a�� �?             =@             
                   =@�LQ�1	�?             7@              	                   �?      �?             @        ������������������������       �                      @        ������������������������       �                      @                              `�b@�}�+r��?             3@       ������������������������       �                     *@                                 �?r�q��?             @       ������������������������       �                     @                                 �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                              ���X@      �?             @        ������������������������       �                     @        ������������������������       �                     @                                 �?      �?             @        ������������������������       �                     @        ������������������������       �                     @                                 �?�����?             3@                                �?�eP*L��?             &@       ������������������������       �                     @                                �K@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �t�bh�h*h-K ��h/��R�(KMKK��h]�B�       �|@     �o@     �y@     �e@      5@      A@       @      ;@      �?      ;@      �?      �?              �?      �?                      :@      �?              3@      @       @      @              @       @              1@      �?      $@              @      �?      @              �?      �?              �?      �?             px@     �a@     �E@      �?      &@              @@      �?      0@              0@      �?      $@              @      �?              �?      @             �u@     `a@     �J@     �X@      @      J@      @      1@      @       @              @      @      @              �?      @       @      @                       @              "@             �A@      I@      G@      >@      G@      =@      B@       @              ;@      B@       @      1@       @      @       @      �?              �?       @                      @              (@      9@      3@      9@      .@      @      "@      @      @      @      @      @      @      @       @               @      @                      @              �?      �?                       @      4@      @      $@      �?      $@                      �?      $@      @      "@      @      @      @      �?      �?              �?      �?              @       @      @                       @      @       @               @      @              �?                      @      �?      $@              $@      �?              4@             pr@     �D@     �B@      &@     �A@      &@      A@      "@      0@      @               @      0@      @               @      0@      @      "@      @      @              @      @      �?      @      @              @              2@       @      $@       @      @              @       @      @      �?      �?      �?      �?                      �?      @                      �?       @              �?       @               @      �?               @              p@      >@              �?      p@      =@      5@       @      5@      @      (@      @      $@      @              �?      $@       @      @              @       @               @      @               @      @              @       @              "@      �?      @              @      �?      �?      �?              �?      �?               @                      �?     �m@      5@      e@      2@     �d@      0@     �B@       @       @             �A@       @      9@       @      (@       @      $@               @       @       @                       @      *@              $@             @`@      ,@      O@      @     �C@      @      *@      �?      $@      �?      @              @      �?      @      �?      �?              @              :@       @      &@              .@       @      &@              @       @              �?      @      �?       @               @      �?              �?       @              7@              Q@      &@     @P@      &@      �?              P@      &@     �F@      &@              @     �F@       @      "@              B@       @      @       @     �@@      @      =@      @      3@              $@      @              �?      $@       @       @      �?       @                      �?       @      �?       @      �?      @              @      @      @              �?      @              @      �?              3@              @               @       @               @       @              Q@      @      .@             �J@      @      $@      @      @      @              @      @              @             �E@             �F@     @T@      C@     @T@      9@     �R@      6@      R@      @      <@              0@      @      (@      �?      "@              @      �?      @               @      �?      �?      �?                      �?       @      @      �?              �?      @      �?                      @      3@      F@      *@      5@      @      @      @       @      �?      �?              �?      �?              @      �?      �?      @              @      �?              @      ,@              (@      @       @       @       @      �?              �?       @      �?                       @      @              @      7@      @      4@       @       @       @                       @      �?      2@              *@      �?      @              @      �?       @               @      �?              @      @              @      @              @      @              @      @              *@      @      @      @              @      @      �?      @                      �?       @              @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJS�)/hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM?huh*h-K ��h/��R�(KM?��h|�B�O         �                    �?�1�uџ�?�           @�@              C                     �?�)85̻�?X           �@               .                 03�I@*;L]n�?M             ^@              -                    �?�z�G��?'             N@              
                    �?�k��(A�?&            �M@                                ���;@r�q��?             @        ������������������������       �                     @               	                   �B@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               ,                 `f�B@�T`�[k�?#            �J@                               ���=@����X�?             E@                                  �?�LQ�1	�?             7@                                ���<@r�q��?             @        ������������������������       �                      @                                  �E@      �?             @        ������������������������       �                     �?        ������������������������       �                     @                                ��$:@�t����?             1@        ������������������������       �                     @                                03k:@r�q��?             (@        ������������������������       �                     �?                                `f�;@�C��2(�?             &@                                  H@ףp=
�?             $@        ������������������������       �                     @                                  @L@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?               +                   �Q@�\��N��?             3@                                   �?j���� �?             1@        ������������������������       �                     @        !       "                   �;@�θ�?
             *@        ������������������������       �                     �?        #       *                   �J@r�q��?	             (@       $       )                   �H@�<ݚ�?             "@       %       &                   �A@      �?              @       ������������������������       �                     @        '       (                   @B@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �                     �?        /       8                   �D@r�q��?&             N@       0       1                    �?�}�+r��?             C@       ������������������������       �                     <@        2       5                    �?z�G�z�?             $@        3       4                 �U�X@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        6       7                 03�P@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        9       <                   �G@���|���?             6@        :       ;                    �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        =       >                    �?�r����?             .@        ������������������������       �                      @        ?       @                 @�pX@8�Z$���?             *@       ������������������������       �                     $@        A       B                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        D       w                    �?f��>���?           �z@        E       n                    =@�ʻ����?=            �Y@       F       ]                    �?� �	��?+            �R@        G       X                   P,@�Gi����?            �B@       H       K                   �5@��X��?             <@        I       J                    3@���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        L       M                   �;@��+7��?             7@        ������������������������       �                     @        N       O                 0��@      �?
             0@        ������������������������       �                     @        P       Q                 ���@      �?             (@        ������������������������       �                     @        R       S                 ���@�q�q�?             "@        ������������������������       �                     @        T       W                 pF @      �?             @       U       V                 �&B@���Q��?             @       ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                     �?        Y       Z                   �6@�q�q�?             "@        ������������������������       �                     @        [       \                 pF�-@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ^       e                     @p9W��S�?             C@        _       b                   �9@�q�q�?             (@       `       a                   �6@r�q��?             @        ������������������������       �                     @        ������������������������       ��q�q�?             @        c       d                 03�0@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        f       g                 ���@8�Z$���?             :@        ������������������������       �                      @        h       i                   �9@�8��8��?             8@       ������������������������       �        	             0@        j       m                    ;@      �?              @        k       l                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        o       p                   @B@�����H�?             ;@       ������������������������       �        
             1@        q       v                    �?�z�G��?             $@       r       s                     @�<ݚ�?             "@       ������������������������       �                     @        t       u                    K@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        x       �                     @��e�1�?�            0t@        y       |                    4@���}<S�?.            @Q@        z       {                    &@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        }       ~                    ?@��S�ۿ?(             N@        ������������������������       �                     @@               �                   �*@؇���X�?             <@        �       �                 ��Y)@���!pc�?	             &@        ������������������������       �                     @        �       �                   @B@      �?             @        ������������������������       �                      @        �       �                   @D@      �?             @        ������������������������       �                     �?        �       �                   �G@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        �       �                    @@�IєX�?             1@        ������������������������       �                     �?        ������������������������       �        
             0@        �       �                  �v6@�i��b��?�            �o@       �       �                   �;@�y)|���?�            @n@        �       �                   �:@b:�&���?7            �T@       �       �                 ��q1@R���Q�?4             T@       �       �                 ��Y @�r����?2            �R@       �       �                    �?�>4և��?%             L@        �       �                   �7@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    1@���c���?"             J@        �       �                 pf�@և���X�?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        �       �                 @3�@��S�ۿ?            �F@       �       �                 ��@г�wY;�?             A@        ������������������������       �                     2@        �       �                 �?$@      �?             0@        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        
             *@        �       �                   �3@"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     3@        �       �                   �2@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                 @3�@ E�+0+�?c            �c@       �       �                    �?�Ι����?:            @X@        �       �                   @@z�G�z�?             9@       �       �                   @<@ףp=
�?             4@       �       �                 ���@"pc�
�?             &@        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     "@        �       �                   �<@���Q��?             @        ������������������������       �                     �?        �       �                    ?@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?      �?+             R@        �       �                    �?�8��8��?             8@       �       �                   �<@�����?             5@       �       �                  s�@�IєX�?
             1@        ������������������������       �                     @        �       �                 ��(@�8��8��?             (@       ������������������������       �؇���X�?             @        ������������������������       �                     @        �       �                    >@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?8��8���?             H@       �       �                 �?�@*
;&���?             G@       �       �                   �@$�q-�?            �C@       �       �                 �&B@؇���X�?             5@       �       �                 ���@ףp=
�?
             4@       ������������������������       �                     *@        �       �                   �>@����X�?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             2@        �       �                   �?@և���X�?             @        ������������������������       �                     �?        �       �                   �D@      �?             @       �       �                   �A@���Q��?             @       ������������������������       ��q�q�?             @        ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    ?@�g�y��?)             O@       �       �                 �̜!@@��8��?             H@        �       �                   �<@���7�?             6@       �       �                 ��) @�X�<ݺ?             2@       ������������������������       �        
             1@        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     :@        �       �                    �?@4և���?             ,@        ������������������������       �                     �?        �       �                   @@@$�q-�?             *@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             &@        �       �                    ;@�8��8��?             (@        ������������������������       �                     @        �       �                    �?�����H�?             "@       �       �                    >@r�q��?             @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     @        �                           @"�!���?q            �d@        �       �                    �?     ��?5             T@        �       �                    �?�t����?             1@       ������������������������       �                     "@        �       �                     �?      �?              @       �       �                   @B@և���X�?             @       �       �                    �?���Q��?             @        ������������������������       �                      @        �       �                    6@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �2@��d��?(            �O@        �       �                     �?���7�?             6@        �       �                 ���`@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     .@        �                       03c@��P���?            �D@       �                       ���`@�c�Α�?             =@              	                   �?�<ݚ�?             ;@                                �=@�q�q�?             "@                               �E@r�q��?             @                               �A@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                                 �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        
                         �?r�q��?             2@       ������������������������       �        	             *@                                  �?���Q��?             @                               @F@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @                              `f�m@�8��8��?             (@       ������������������������       �                     "@                                 �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?              *                   �?>���Rp�?<            �U@                              P��%@r�q��?             8@                              �(\�?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @              )                   �?�q�q�?             2@             (                   @      �?             0@             %                   �?����X�?             ,@              $                ���.@�q�q�?             @              #                   �?�q�q�?             @       !      "                P��+@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        &      '                `f7@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        +      8                   @�? Da�?+            �O@       ,      -                   @     ��?             @@        ������������������������       �                     @        .      3                   �?�>����?             ;@        /      2                  �<@ףp=
�?             $@        0      1                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        4      7                   �?�IєX�?             1@        5      6                  �1@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             *@        9      >                ���A@�g�y��?             ?@        :      ;                ��T?@$�q-�?	             *@       ������������������������       �                     &@        <      =                   @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     2@        �t�bh�h*h-K ��h/��R�(KM?KK��h]�B�       P|@     0p@     @w@     �e@      J@      Q@      E@      2@      E@      1@      �?      @              @      �?      �?              �?      �?             �D@      (@      >@      (@      4@      @      @      �?       @              @      �?              �?      @              .@       @      @              $@       @              �?      $@      �?      "@      �?      @              @      �?              �?      @              �?              $@      "@      $@      @              @      $@      @              �?      $@       @      @       @      @      �?      @              �?      �?              �?      �?                      �?      @                       @      &@                      �?      $@      I@       @      B@              <@       @       @      �?      @              @      �?              �?      @              @      �?               @      ,@      @      �?              �?      @               @      *@               @       @      &@              $@       @      �?       @                      �?      t@     @Z@     �F@     �L@      E@     �@@      .@      6@      "@      3@      @       @               @      @              @      1@              @      @      $@              @      @      @      @              @      @              @      @      @       @      @       @       @              �?      �?              @      @      @              �?      @      �?                      @      ;@      &@      @      @      �?      @              @      �?       @      @       @               @      @              6@      @               @      6@       @      0@              @       @      @       @               @      @              @              @      8@              1@      @      @       @      @              @       @       @       @                       @      �?             0q@      H@     �O@      @      @       @               @      @              L@      @      @@              8@      @       @      @      @              @      @               @      @      �?      �?               @      �?      �?      �?      �?              0@      �?              �?      0@             �j@      E@     `j@      ?@      Q@      .@      Q@      (@     @P@      $@      G@      $@      �?      @              @      �?             �F@      @      @      @      �?               @      @      E@      @     �@@      �?      2@              .@      �?       @      �?       @                      �?      *@              "@       @               @      "@              3@              @       @      @                       @              @     �a@      0@     �T@      ,@      4@      @      2@       @      "@       @      @              @       @      "@               @      @      �?              �?      @              @      �?             �O@      "@      6@       @      3@       @      0@      �?      @              &@      �?      @      �?      @              @      �?              �?      @              @             �D@      @     �C@      @      B@      @      2@      @      2@       @      *@              @       @      @       @      �?                      �?      2@              @      @              �?      @      @      @       @       @      �?      �?      �?              �?       @              N@       @     �G@      �?      5@      �?      1@      �?      1@                      �?      @              :@              *@      �?      �?              (@      �?      �?      �?              �?      �?              &@              �?      &@              @      �?       @      �?      @      �?       @              @              @     @T@     �U@      .@     @P@      @      (@              "@      @      @      @      @       @      @               @       @      �?              �?       @               @              �?              $@     �J@      �?      5@      �?      @              @      �?                      .@      "@      @@       @      5@      @      5@      @      @      �?      @      �?       @               @      �?                      @       @      �?              �?       @              @      .@              *@      @       @      �?       @               @      �?               @               @              �?      &@              "@      �?       @               @      �?             �P@      5@      &@      *@      @      �?              �?      @              @      (@      @      (@      @      $@       @      @       @      �?      �?      �?              �?      �?              �?                      @       @      @              @       @                       @       @             �K@       @      9@      @              @      9@       @      "@      �?      �?      �?              �?      �?               @              0@      �?      @      �?      @                      �?      *@              >@      �?      (@      �?      &@              �?      �?              �?      �?              2@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ[س=hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM1huh*h-K ��h/��R�(KM1��h|�B@L         \                    �?l��n�?�           @�@                                    @��'�e��?�            `l@                                  @�-���e�?N            �_@        ������������������������       �                      @                                   �?Ȓ�g;�?M             _@                                0Cd=@������?             B@               
                    �?؇���X�?             @              	                 03[:@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     =@                                   �?�C��2(�?3             V@                                   �?$�q-�?,            �S@        ������������������������       �                     <@                                   �?H%u��?             I@                                  6@(L���?            �E@                                  �?d}h���?             <@                               `f�)@8�Z$���?             :@        ������������������������       �                     @                                   :@z�G�z�?	             4@        ������������������������       �և���X�?             @        ������������������������       �                     *@        ������������������������       �                      @        ������������������������       �        	             .@        ������������������������       �                     @                                ���[@z�G�z�?             $@       ������������������������       �                     @                                  �8@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                I                    �?&�����?C            @Y@       !       D                  S�-@�ɞ`s�?*            �N@       "       -                 ��@8�A�0��?              F@        #       $                 03�@���N8�?             5@        ������������������������       �                     �?        %       ,                    �?z�G�z�?             4@       &       '                    �?�S����?             3@        ������������������������       �                     @        (       )                   �5@z�G�z�?
             .@        ������������������������       �                      @        *       +                 ���@$�q-�?	             *@        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                     �?        .       /                    �?\X��t�?             7@        ������������������������       �                      @        0       1                    �?�G��l��?             5@        ������������������������       �                      @        2       A                   �=@D�n�3�?             3@       3       4                    0@�	j*D�?
             *@        ������������������������       �                      @        5       >                 @�"@���|���?	             &@       6       =                    ;@      �?              @       7       <                   �9@�q�q�?             @       8       ;                   �7@z�G�z�?             @        9       :                    5@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ?       @                 �[$@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        B       C                    A@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        E       F                 03�1@�IєX�?
             1@       ������������������������       �                     *@        G       H                    7@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        J       U                    �?H�z�G�?             D@        K       T                 `f7@      �?
             0@       L       M                    @؇���X�?	             ,@        ������������������������       �                     �?        N       S                    �?$�q-�?             *@        O       P                    �?z�G�z�?             @        ������������������������       �                     @        Q       R                   �<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        V       [                    @�q�q�?             8@        W       X                    @r�q��?             @        ������������������������       �                     @        Y       Z                    @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     2@        ]       d                    @��.D��?0           P~@        ^       _                    @�4�����?             ?@       ������������������������       �                     3@        `       a                 ��T?@r�q��?             (@       ������������������������       �                     @        b       c                 ���A@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        e       �                     �?�X��M�?           `|@        f       �                 @�:x@��J���?@            �Z@       g       �                 �D�M@�B�����?>             Z@       h       q                    �?h+�v:�?)             Q@        i       j                   �:@      �?             (@        ������������������������       �                     @        k       p                    �?�q�q�?             "@       l       m                 ���<@      �?              @        ������������������������       �                     @        n       o                   �B@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        r       s                 ��$:@X�Cc�?"             L@        ������������������������       �                     @        t       �                    �?���Q��?             I@       u       |                   �@@\�Uo��?             C@        v       {                   �<@@4և���?             ,@       w       z                 `f�D@�C��2(�?             &@        x       y                   �@@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        }       �                   �J@�q�q�?             8@       ~       �                 �T!@@������?
             1@              �                   `G@�r����?             .@       �       �                 `f�;@����X�?             @       �       �                   �E@r�q��?             @        ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                 `fF<@؇���X�?             @        ������������������������       �                     @        �       �                   @>@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�q�q�?             (@       �       �                 `fFJ@�z�G��?             $@        ������������������������       �                     @        �       �                   @D@      �?             @       �       �                    7@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?4?,R��?             B@       �       �                   �G@����X�?             ,@       �       �                    �?      �?              @       �       �                   �;@r�q��?             @        �       �                   �8@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?      �?             @       �       �                 @�pX@���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?���7�?
             6@        �       �                 `��W@�8��8��?             (@        �       �                    �?z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                     @        �       *                �T�I@���3���?�            �u@       �       )                   �?dk�����?�             u@       �       �                    �?������?�            t@        �       �                   @@dP-���?            �G@        ������������������������       �                     9@        �       �                    �?"pc�
�?             6@       �       �                   �8@d}h���?	             ,@        ������������������������       �                     @        �       �                 ��%@���!pc�?             &@       �       �                   �<@      �?              @        ������������������������       �                     @        �       �                    ?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ���,@�q�q�?             @        ������������������������       �                     �?        �       �                    ;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ��3@      �?              @        �       �                    7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       $                   �?��cd@�?�             q@       �                         @@@�G�c��?�            �o@       �       �                 ���@p*aƿ �?|             h@        �       �                 `f�@      �?             (@       �       �                     @      �?              @        ������������������������       �                      @        �       �                    6@      �?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                    :@      �?             @       �       �                 �&b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                  ��@��/�8�?u            �f@        ������������������������       �                     6@        �                         �?@�W��}�?i            �c@       �                       ���#@h������?d            �b@       �       �                   �<@�϶O'3�?G            @Z@       �       �                    �?�9�a��?@            �W@       �       �                   �0@��{H�?:            �U@        ������������������������       �      �?              @        �       �                 ��) @,�"���?8            @U@       �       �                 �1@ ����?-            @P@        �       �                 ��@"pc�
�?             6@        �       �                    7@�C��2(�?             &@        ������������������������       �                     @        ������������������������       �      �?              @        �       �                   �3@���!pc�?             &@        ������������������������       �                      @        �       �                 �?$@�q�q�?             "@        �       �                    ;@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        �       �                   �5@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �?�@Du9iH��?            �E@       ������������������������       �                     7@        �       �                   �4@R���Q�?             4@        ������������������������       �      �?             @        ������������������������       �                     0@        �       �                   �9@�z�G��?             4@       ������������������������       �                     &@        �       �                 pf� @�q�q�?             "@        ������������������������       �                     @        �       �                 ��)"@      �?             @       �       �                   �;@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?և���X�?             @        ������������������������       �                     �?        �       �                   �9@      �?             @        ������������������������       �                     @        ������������������������       �                     @        �                          �=@�eP*L��?             &@       �       �                    �?����X�?             @        ������������������������       �                     @        �       �                 ���"@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @                                 ;@���.�6�?             G@        ������������������������       �                     4@                                 �?ȵHPS!�?             :@             
                    @ �q�q�?             8@              	                   �?�8��8��?             (@                               �<@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                      @                              ��i @      �?              @        ������������������������       �                     @                                  @z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @                              �?�@�g�y��?+             O@        ������������������������       �                     8@                                  @�}�+r��?             C@                               �*@���7�?             6@                             `f�)@@4և���?             ,@       ������������������������       �                     @                                @D@؇���X�?             @        ������������������������       �                     @                                 G@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @              #                @3�@      �?             0@              "                   �?z�G�z�?             @              !                  �D@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     &@        %      &                  x@@�KM�]�?             3@       ������������������������       �        	             (@        '      (                   @����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        	             .@        +      0                   >@���|���?             &@       ,      /                   ;@և���X�?             @       -      .                   6@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �t�b�      h�h*h-K ��h/��R�(KM1KK��h]�B       {@     pq@     �J@     �e@      &@     �\@       @              "@     �\@      �?     �A@      �?      @      �?      @              @      �?                       @              =@       @      T@      @      R@              <@      @      F@      @     �B@      @      6@      @      6@              @      @      0@      @      @              *@       @                      .@              @       @       @              @       @      �?              �?       @              E@     �M@      3@      E@      2@      :@      @      0@      �?              @      0@      @      0@              @      @      (@       @              �?      (@      �?                      (@      �?              *@      $@       @              &@      $@               @      &@       @      "@      @       @              @      @      @       @      @       @      @      �?      �?      �?      �?                      �?      @                      �?       @              �?       @               @      �?               @      @              @       @              �?      0@              *@      �?      @      �?                      @      7@      1@      @      (@       @      (@      �?              �?      (@      �?      @              @      �?      �?      �?                      �?               @       @              3@      @      �?      @              @      �?       @      �?                       @      2@             �w@     @Z@      $@      5@              3@      $@       @      @              @       @               @      @              w@      U@     @R@      A@     @R@      ?@      E@      :@      @      @              @      @      @      @      @      @              �?      @              @      �?              �?              B@      4@      @              >@      4@      7@      .@      *@      �?      $@      �?      @      �?      @                      �?      @              @              $@      ,@      @      *@       @      *@       @      @      �?      @              @      �?       @      �?                       @       @              @      �?      @              @      �?              �?      @              @      @      @      @      @              @      @      �?      @      �?                      @       @                       @      ?@      @      $@      @      @      �?      @      �?       @      �?       @                      �?      @               @              @      @      @       @               @      @                      �?      5@      �?      &@      �?      @      �?      @                      �?      @              $@                      @     �r@      I@     Pr@     �E@     `q@     �E@     �E@      @      9@              2@      @      &@      @      @               @      @      @      �?      @               @      �?              �?       @              �?       @              �?      �?      �?              �?      �?              @      �?       @      �?              �?       @              @             `m@     �C@     @k@     �B@     �c@     �A@      @      @      @      @       @              @      @      @                      @      �?      @      �?      �?      �?                      �?               @      c@      =@      6@             @`@      =@     �_@      9@     �T@      6@     @S@      1@     @R@      ,@      �?      �?      R@      *@      M@      @      2@      @      $@      �?      @              @      �?       @      @       @              @      @       @       @      �?              �?       @      @      �?              �?      @              D@      @      7@              1@      @      �?      @      0@              ,@      @      &@              @      @              @      @      @       @      @              @       @              �?              @      @      �?              @      @              @      @              @      @       @      @              @       @       @       @                       @      @             �E@      @      4@              7@      @      7@      �?      &@      �?      $@      �?              �?      $@              �?              (@                       @      @      @              @      @      �?              �?      @              N@       @      8@              B@       @      5@      �?      *@      �?      @              @      �?      @              @      �?              �?      @               @              .@      �?      @      �?       @      �?       @                      �?       @              &@              1@       @      (@              @       @               @      @              .@              @      @      @      @      �?      @      �?                      @      @                      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJnխphG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM%huh*h-K ��h/��R�(KM%��h|�B@I         Z                    �?z��Y�)�?�           @�@               Y                    @~�1u���?�            @k@              N                    @���N8�?�            @j@              G                    @@�'�`d�?~            �h@                                   @��c����?X             a@                                   �?ףp=
�?%             N@        ������������������������       �                     5@                                   �?8�Z$���?            �C@       	                           6@     ��?             @@        
                           �?���Q��?             @                                  :@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     ;@                                ���`@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @               :                    �?�eP*L��?3            @S@                                  �?�w��#��?#             I@                                H�%@�����H�?             "@       ������������������������       �                     @                                   �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @               7                    �?hP�vCu�?            �D@              &                    �?؀�:M�?            �B@                                   1@�t����?
             1@        ������������������������       �                     @                                �&�@�q�q�?             (@        ������������������������       �                      @                !                    9@�z�G��?             $@        ������������������������       �                      @        "       %                 pF @      �?              @       #       $                 �&B@r�q��?             @       ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        '       ,                 @3�@�G�z��?             4@        (       )                 P��@z�G�z�?             $@        ������������������������       �                     @        *       +                   �9@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        -       6                 ��&@�z�G��?             $@       .       /                 ��� @�<ݚ�?             "@        ������������������������       �                     @        0       5                   �;@�q�q�?             @       1       4                    4@z�G�z�?             @        2       3                   �#@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        8       9                   �;@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ;       F                 ��Z5@�q�q�?             ;@       <       =                    @և���X�?             5@        ������������������������       �                     @        >       ?                    ;@      �?
             0@        ������������������������       �                     @        @       A                    �?X�<ݚ�?             "@        ������������������������       �                      @        B       C                   �.@����X�?             @        ������������������������       �                     @        D       E                   �=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        H       I                     @��v$���?&            �N@       ������������������������       �        #            �K@        J       K                 `f(@r�q��?             @        ������������������������       �                     @        L       M                   `1@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        O       X                 ���d@�q�q�?
             (@       P       Q                    �?z�G�z�?             $@        ������������������������       �                      @        R       S                 ���1@      �?              @        ������������������������       �                     �?        T       W                     @؇���X�?             @        U       V                 ��T?@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        [       �                    �?X���?�?2           �~@        \       m                   �;@҄��?.            �P@        ]       l                  ��^@�q�q�?             5@       ^       _                     �?�z�G��?             4@        ������������������������       �                     @        `       a                    @և���X�?
             ,@        ������������������������       �                     @        b       c                     @�q�q�?             "@        ������������������������       �                      @        d       g                 ���@և���X�?             @        e       f                   �7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        h       i                 �0@      �?             @        ������������������������       �                      @        j       k                   �2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        n       y                     �?z�G�z�?             �F@        o       x                 @�ys@�E��ӭ�?             2@       p       u                    �?     ��?             0@       q       t                 `f�B@8�Z$���?	             *@       r       s                 ��>@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        v       w                   �K@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        z       �                   �=@PN��T'�?             ;@       {       �                 H�Z&@z�G�z�?             4@       |       �                   @@      �?
             0@       }       ~                 ���@8�Z$���?             *@        ������������������������       �                      @               �                   @<@"pc�
�?             &@       ������������������������       �z�G�z�?             $@        ������������������������       �                     �?        �       �                   �<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    @T�����?           �z@        �       �                     @������?             .@        ������������������������       �                     @        �       �                     @      �?              @        ������������������������       �                     @        �       �                    �?z�G�z�?             @       ������������������������       �                     @        �       �                 ��T?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �                         �C@(2��R�?�            �y@       �                          @��Ex�?�            Pt@       �                          �?ihh��?�            ps@       �       �                 ��D:@�;n��?�            @s@       �       �                 ��i @��-���?�            p@       �       �                 ��) @.�w��K�?]            �b@       �       �                    �?��
CJ�?\            `b@        �       �                    �?�C��2(�?             6@       �       �                  s�@�����?             5@        ������������������������       �                      @        �       �                   �=@8�Z$���?             *@       ������������������������       �z�G�z�?             $@        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�J�4�?N            @_@       �       �                    �?�<�}���?L            @^@       �       �                   �;@r�q��?K             ^@        �       �                    �? {��e�?#            �J@       �       �                 ��@&^�)b�?            �E@        ������������������������       �                     @        �       �                   �5@�˹�m��?             C@        �       �                 @3�@��2(&�?             6@       �       �                   �4@      �?
             0@       ������������������������       �                     "@        �       �                 ��L@؇���X�?             @        �       �                  s@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �1@�q�q�?             @        ������������������������       �                     �?        �       �                   �3@���Q��?             @       ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                     0@        �       �                 P�@�z�G��?             $@       �       �                   �7@      �?              @        ������������������������       �                     @        �       �                   �9@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                     @��v����?(            �P@        ������������������������       �                     *@        �       �                 @3�@r�q��?"             K@       �       �                 �?�@�<ݚ�?             B@       �       �                 �?$@H%u��?             9@        �       �                    =@���!pc�?             &@       �       �                 pf�@�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     ,@        �       �                   �?@�eP*L��?             &@        ������������������������       �                      @        �       �                   �A@�q�q�?             "@       ������������������������       �z�G�z�?             @        ������������������������       �      �?             @        �       �                    ?@�X�<ݺ?
             2@       ������������������������       �                     .@        �       �                   �@@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                 03�6@�8��8��?@             [@       �       �                   �<@�8��8N�?5             X@       �       �                   �*@����1�?*            @R@       �       �                     @L紂P�?            �I@        �       �                   �(@���N8�?             5@        �       �                   �2@z�G�z�?             @        ������������������������       �                      @        �       �                   �5@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �;@      �?             0@       ������������������������       �                     (@        ������������������������       �                     @        �       �                 ���!@��S�ۿ?             >@        �       �                 pf� @؇���X�?             ,@        ������������������������       �                      @        �       �                    �?r�q��?             (@       �       �                    8@"pc�
�?             &@       ������������������������       �                     @        �       �                   �;@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             0@        ������������������������       �                     6@        ������������������������       �                     7@        �       �                    �?r�q��?             (@       �       �                   �@@"pc�
�?
             &@       �       �                 03�7@����X�?             @        ������������������������       �                     �?        �       �                    >@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �                          �?ҳ�wY;�?            �I@       �                          �?�û��|�?             G@       �                         �?@�q�q�?             B@       �       �                   �>@�z�G��?             >@        �       �                   @>@�<ݚ�?             "@       �       �                   �<@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �                           7@�����?             5@        ������������������������       �                     @                              0�K@�����H�?
             2@                             ��yC@@4և���?             ,@                                �@@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �      �?             @        ������������������������       �                     @        	                      03U@�z�G��?             $@       
                      ���M@      �?              @                                =@      �?             @                                7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @                                   @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        
             ,@                                 �?�zvܰ?0             V@        ������������������������       �                     &@              "                   �?`<)�+�?,            @S@             !                   �?��
���?*            �R@                               @I@�]0��<�?#            �N@        ������������������������       �                     A@                              `fF:@�>����?             ;@       ������������������������       �        
             0@                                 @J@"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     ,@        #      $                     @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �t�bh�h*h-K ��h/��R�(KM%KK��h]�BP       �|@     @o@      M@      d@      I@      d@      E@     �c@     �D@      X@      @      K@              5@      @     �@@      @      =@      @       @       @       @       @                       @      �?                      ;@      @      @              @      @             �A@      E@      1@     �@@      �?       @              @      �?      @      �?                      @      0@      9@      ,@      7@      @      (@              @      @      @       @              @      @               @      @      @      �?      @      �?       @              @       @              "@      &@       @       @              @       @      @       @                      @      @      @      @       @      @              @       @      @      �?      �?      �?              �?      �?              @                      �?              �?       @       @               @       @              2@      "@      (@      "@              @      (@      @      @              @      @               @      @       @      @              �?       @               @      �?              @              �?      N@             �K@      �?      @              @      �?       @      �?                       @       @      @       @       @       @              @       @              �?      @      �?       @      �?       @                      �?      @                       @       @             @y@     �V@     �E@      7@      @      ,@      @      ,@              @      @       @              @      @      @       @              @      @      �?       @               @      �?              @      �?       @              �?      �?      �?                      �?      �?              B@      "@      *@      @      *@      @      &@       @      @       @      @                       @      @               @      �?       @                      �?               @      7@      @      0@      @      (@      @      &@       @       @              "@       @       @       @      �?              �?       @      �?                       @      @              @             �v@     �P@      @      &@              @      @      @              @      @      �?      @              �?      �?      �?                      �?     Pv@      L@      q@     �J@      p@     �J@     p@     �I@      l@     �@@     @_@      8@     @_@      6@      4@       @      3@       @       @              &@       @       @       @      @              �?             @Z@      4@     @Y@      4@      Y@      4@      E@      &@     �A@       @              @     �A@      @      3@      @      .@      �?      "@              @      �?      �?      �?      �?                      �?      @              @       @      �?              @       @       @       @      �?              0@              @      @      @      �?      @              @      �?              �?      @                       @      M@      "@      *@             �F@      "@      <@       @      6@      @       @      @      @      @      @                      @       @              ,@              @      @               @      @      @      @      �?       @       @      1@      �?      .@               @      �?              �?       @              �?              @                       @     �X@      "@     @V@      @     �P@      @      F@      @      0@      @      @      �?       @               @      �?              �?       @              (@      @      (@                      @      <@       @      (@       @       @              $@       @      "@       @      @              @       @               @      @              �?              0@              6@              7@              $@       @      "@       @      @       @              �?      @      �?      @                      �?      @              �?             �@@      2@      <@      2@      5@      .@      5@      "@       @      @       @      @              @       @                      @      3@       @      @              0@       @      *@      �?      @      �?      @                      �?      "@              @      �?              @      @      @      @      �?      @      �?      �?      �?      �?                      �?       @              @                       @      @              �?       @               @      �?              ,@             @U@      @      &@             �R@      @     @R@       @     �M@       @      A@              9@       @      0@              "@       @               @      "@              ,@              �?      �?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�[�.hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM/huh*h-K ��h/��R�(KM/��h|�B�K         d                    �?@?�p�?�           @�@               _                 p�H@�+��0��?�             p@              &                 `f�$@      �?s             h@               %                    �?~|z����?"            �J@                                  -@�q���?             H@        ������������������������       �                     @               $                    �?X�<ݚ�?            �F@              	                    1@�eP*L��?             F@        ������������������������       �                     @        
       #                    K@�p ��?            �D@                               ���@Hث3���?            �C@                                   �?؇���X�?             ,@                               �Y�@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @                                �̌@ �o_��?             9@                                  �?��
ц��?	             *@                               �&B@և���X�?             @                                 �5@      �?             @        ������������������������       �                      @                                   9@      �?             @        ������������������������       �                      @        ������������������������       �      �?              @        ������������������������       �                     �?                                   4@�q�q�?             @        ������������������������       �                     @                                ��@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @               "                   �;@�8��8��?             (@                !                    9@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        '       X                    @2�ߣ0��?Q            `a@       (       W                    @d58��1�?J            �^@       )       >                    �?R���Q�?H             ^@       *       1                     @؇���X�?&             L@       +       0                    �?P���Q�?             D@       ,       /                    �? 	��p�?             =@        -       .                 `v7<@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     8@        ������������������������       �                     &@        2       7                    �?      �?             0@        3       4                 ��&@�q�q�?             @        ������������������������       �                     �?        5       6                 ���*@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        8       =                 �A7@�	j*D�?             *@       9       <                    �?"pc�
�?             &@        :       ;                 ��*@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ?       J                    �?     ��?"             P@        @       A                   �,@ �Cc}�?             <@        ������������������������       �                     @        B       C                     @؇���X�?             5@        ������������������������       �                     @        D       E                   @5@d}h���?             ,@        ������������������������       �                     �?        F       I                    �?8�Z$���?             *@        G       H                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        K       L                     @X�<ݚ�?             B@        ������������������������       �                     .@        M       N                    @���N8�?             5@        ������������������������       �                      @        O       V                 ��1@�S����?
             3@        P       U                    �?և���X�?             @       Q       R                 @3�/@      �?             @        ������������������������       �                     �?        S       T                    ;@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                      @        Y       Z                    @�t����?             1@        ������������������������       �                     @        [       \                 ��T?@z�G�z�?             $@        ������������������������       �                     @        ]       ^                    %@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        `       c                     @�FVQ&�?(            �P@       a       b                     @      �?&             P@        ������������������������       �                      @        ������������������������       �        %             O@        ������������������������       �                      @        e       �                    �?>.��Y��?*           `|@        f       }                     �?8����?/            @Q@        g       t                    �?�f7�z�?             =@       h       s                   �A@�ՙ/�?             5@       i       j                 ���<@��S���?             .@        ������������������������       �                     @        k       p                  "&d@�q�q�?             (@       l       m                 `f�A@؇���X�?             @        ������������������������       �                     @        n       o                 �M@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        q       r                 p�w@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        u       v                 ��+T@      �?              @        ������������������������       �                     @        w       x                 ��hU@z�G�z�?             @        ������������������������       �                      @        y       |                    �?�q�q�?             @       z       {                 p"�X@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ~       �                    5@R���Q�?             D@               �                 ؼC1@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �=@؇���X�?            �A@       �       �                   �<@��<b���?             7@       �       �                    �?؇���X�?             5@       �       �                 83�0@R���Q�?             4@       �       �                   @@�����H�?             2@       �       �                 ���@z�G�z�?	             $@        ������������������������       �                     @        �       �                    9@����X�?             @        ������������������������       �                     �?        �       �                   @<@�q�q�?             @       ������������������������       ����Q��?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     (@        �       �                     �?z���=��?�            x@        �       �                 ��yC@�q�q�?)            �P@       �       �                   �9@��Zy�?            �C@        ������������������������       �                     @        �       �                 03k:@     ��?             @@        ������������������������       �                      @        �       �                   �J@      �?             >@       �       �                   �;@�q�q�?             5@        ������������������������       �                      @        �       �                 `f�;@p�ݯ��?
             3@        ������������������������       �                     @        �       �                   @>@��S���?             .@        ������������������������       �                      @        �       �                   �>@�n_Y�K�?             *@        ������������������������       �                     @        �       �                   @B@X�<ݚ�?             "@       �       �                   �A@      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    R@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        �       �                    '@�+$�jP�?             ;@        ������������������������       �                     @        �       �                   �B@�8��8��?             8@        �       �                    �?r�q��?             (@       �       �                    >@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             (@        �       .                   @X�(7��?�            �s@       �       %                   B@Pl֕���?�            �r@       �                          �?$�`��S�?�            �q@       �                          �?ܔQ|ӭ�?�            �k@       �                         �N@�:	p��?�            `j@       �                         �C@ ���g=�?�            �i@       �       
                  �*@4�<����?}            @f@       �       �                    �?*.>h�<�?r             d@        �       �                  ��@��s����?             5@        ������������������������       �                     @        �       �                   �<@������?
             .@       �       �                 ��(@"pc�
�?             &@       ������������������������       �z�G�z�?             $@        ������������������������       �                     �?        �       �                    >@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                 03s@؇���X�?c            �a@        �       �                 `f�@�	j*D�?             *@       �       �                     @"pc�
�?             &@       ������������������������       �                     @        �       �                    6@�q�q�?             @        ������������������������       �                      @        �       �                   �>@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �                       `fF)@ ��P0�?[            �_@       �       �                     @�KM�]�?R            �\@        ������������������������       �                      @        �       �                 �?$@���C��?K            �Z@        ������������������������       �                     4@        �       �                 �1@(L���??            �U@        �       �                   �8@���Q��?             @       �       �                   �5@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                 �?�@�����H�?<            @T@        �       �                   �@ ��WV�?             :@        �       �                   �:@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     6@        �                         �B@t�6Z���?)            �K@       �       �                 @3�@H�ՠ&��?(             K@        �       �                    :@�q�q�?             @        ������������������������       �                     �?        �       �                   �?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ���!@�t����?%            �I@       �       �                 pf� @�ݜ�?            �C@       �       �                    4@<���D�?            �@@        �       �                    1@      �?             @        ������������������������       �                     �?        �       �                   �2@���Q��?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        �       �                    ?@ 7���B�?             ;@       ������������������������       �                     6@        �       �                   �@@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    8@r�q��?             @       ������������������������       �                     @        �       �                   �;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 �y�"@�8��8��?	             (@        ������������������������       �                      @        �                       ���#@ףp=
�?             $@       �       �                   �<@�����H�?             "@       ������������������������       �                     @        �                           ?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?              	                   @@�	j*D�?	             *@                               �:@"pc�
�?             &@       ������������������������       �                     @                                 =@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     1@        ������������������������       �                     =@                                 Q@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     "@              "                   �?     ��?'             P@                                #@�rF���?"            �K@        ������������������������       �                      @                                 5@dP-���?            �G@                              03#,@      �?              @                                3@���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @              !                   �? ���J��?            �C@                             039@ ��WV�?             :@       ������������������������       �        	             0@                                 �@@ףp=
�?             $@                                �<@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             *@        #      $                   �?�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        &      -                ��?P@�	j*D�?             *@       '      *                   �?�q�q�?             @       (      )                   >@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        +      ,                  �>@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     6@        �t�bh�h*h-K ��h/��R�(KM/KK��h]�B�       �{@     �p@      S@     �f@      R@      ^@      <@      9@      7@      9@      @              4@      9@      4@      8@              @      4@      5@      4@      3@       @      (@       @      @       @                      @               @      2@      @      @      @      @      @      @      @       @              �?      @               @      �?      �?              �?      @       @      @              �?       @      �?                       @      &@      �?      @      �?      @                      �?       @                       @              �?      @              F@     �W@      =@     @W@      ;@     @W@       @      H@       @      C@       @      ;@       @      @              @       @                      8@              &@      @      $@       @      �?      �?              �?      �?              �?      �?              @      "@       @      "@       @      @              @       @                      @       @              3@     �F@      @      9@              @      @      2@              @      @      &@      �?               @      &@       @      �?       @                      �?              $@      0@      4@              .@      0@      @               @      0@      @      @      @      @      @              �?      @       @      @                       @      �?              (@               @              .@       @      @               @       @      @              @       @               @      @              @      O@       @      O@       @                      O@       @              w@     �U@      H@      5@      1@      (@      *@       @      @       @      @              @       @      �?      @              @      �?      @      �?                      @      @       @      @                       @      @              @      @              @      @      �?       @               @      �?      �?      �?              �?      �?              �?              ?@      "@      �?      @              @      �?              >@      @      2@      @      2@      @      1@      @      0@       @       @       @      @              @       @      �?              @       @      @       @      �?               @              �?      �?              �?      �?              �?                       @      (@              t@     @P@      F@      6@      6@      1@      @              .@      1@               @      .@      .@      @      ,@               @      @      (@              @      @       @       @              @       @              @      @      @      @      @      @                      @      �?               @      �?       @                      �?      6@      @              @      6@       @      $@       @      $@      �?      $@                      �?              �?      (@             @q@     �E@     �o@     �E@     �n@     �C@     @h@      :@      g@      :@     �f@      8@     @c@      8@      a@      8@      1@      @      @              &@      @      "@       @       @       @      �?               @       @               @       @              ^@      4@      "@      @      "@       @      @              @       @       @               @       @               @       @                       @     �[@      0@     �Y@      (@       @             �W@      (@      4@             �R@      (@       @      @       @      �?              �?       @                       @      R@      "@      9@      �?      @      �?      @                      �?      6@             �G@       @     �G@      @       @      �?      �?              �?      �?              �?      �?             �F@      @      A@      @      =@      @      @      @              �?      @       @       @              �?       @      :@      �?      6@              @      �?              �?      @              @      �?      @              �?      �?              �?      �?              &@      �?       @              "@      �?       @      �?      @               @      �?              �?       @              �?                      �?      "@      @      "@       @      @              @       @               @      @                       @      1@              =@               @       @               @       @              "@             �I@      *@     �E@      (@               @     �E@      @      @      @       @      @       @                      @      @              C@      �?      9@      �?      0@              "@      �?       @      �?       @                      �?      @              *@               @      �?              �?       @              "@      @       @      @      �?       @      �?      �?              �?      �?       @               @      �?              @              6@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ��=hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM%huh*h-K ��h/��R�(KM%��h|�B@I         ~                     @�)�>_M�?�           @�@                                  �'@`՟�G��?�            `s@                                   �?<���D�?            �@@        ������������������������       �                      @                                   �?`Jj��?             ?@                                   �?��S�ۿ?             >@        ������������������������       �                     @                                  �H@�8��8��?             8@       	       
                    @�nkK�?             7@        ������������������������       �                     @                                   &@      �?             0@                                 �5@@4և���?	             ,@                                  �1@r�q��?             @        ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?               y                    �?d'����?�            Pq@              &                    �?\X��t�?�            �o@                                   �?����q�?A            @[@                                 �*@�k~X��?+             R@                                   �?`2U0*��?             9@        ������������������������       �                     @                                   :@�X�<ݺ?             2@        ������������������������       �      �?              @        ������������������������       �                     0@        ������������������������       �                     �G@                                    �?�?�|�?            �B@       ������������������������       �                     6@                !                    �?��S�ۿ?	             .@        ������������������������       �                     @        "       #                   �9@�8��8��?             (@        ������������������������       �                     @        $       %                    <@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        '       6                    ,@      �?X             b@        (       )                    �?ܷ��?��?             =@        ������������������������       �                     �?        *       +                 `f�)@ �Cc}�?             <@        ������������������������       �                      @        ,       5                   �*@ȵHPS!�?             :@       -       .                   �:@H%u��?             9@        ������������������������       �                     $@        /       0                    =@z�G�z�?             .@        ������������������������       �                      @        1       2                    C@$�q-�?             *@       ������������������������       �                      @        3       4                   �F@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        7       8                   �-@��.۽0�?E            �\@        ������������������������       �                      @        9       :                    (@
�ۓQ{�?D            @\@        ������������������������       �                      @        ;       x                    �?���{��??            @Z@       <       w                   �R@r�{o43�?>            �Y@       =       b                    �?��[�8��?=            �Y@       >       C                   �;@ {��e�?#            �J@        ?       B                    �?և���X�?             @       @       A                     �?      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        D       a                    �?�㙢�c�?             G@       E       `                 `f�B@z�G�z�?             D@       F       M                    �?�	j*D�?             :@        G       H                 ���<@      �?             @        ������������������������       �                     �?        I       L                 ��L@@�q�q�?             @       J       K                   �E@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        N       _                     �?���!pc�?             6@       O       ^                   �J@�z�G��?             4@       P       ]                   �H@���Q��?             .@       Q       Z                   �A@X�Cc�?
             ,@       R       Y                   �>@���!pc�?             &@       S       X                    G@      �?             @       T       W                   @B@���Q��?             @       U       V                 `fF<@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        [       \                   @B@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     ,@        ������������������������       �                     @        c       d                    6@���c�H�?            �H@        ������������������������       �                     @        e       v                     �?�%^�?            �E@       f       q                   �H@� �	��?             9@       g       p                    �?�	j*D�?             *@       h       o                 03�U@���|���?             &@       i       j                   �;@�q�q�?             @        ������������������������       �                     �?        k       n                    �?z�G�z�?             @        l       m                    C@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        r       s                    L@r�q��?             (@       ������������������������       �                      @        t       u                 `f�R@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        
             2@        ������������������������       �                     �?        ������������������������       �                      @        z       {                 ���i@ �q�q�?             8@       ������������������������       �                     3@        |       }                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?               �                    �?!��)��?�             y@        �       �                    @�'�=z��?F            �`@       �       �                   �7@������?B            �_@        �       �                    @���!pc�?            �K@        �       �                    @��S���?             .@       �       �                    �?z�G�z�?             $@        ������������������������       �                      @        �       �                   �&@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    )@z�G�z�?             D@        ������������������������       �                     &@        �       �                    �?>���Rp�?             =@       �       �                 �[$@ �o_��?             9@       �       �                   �0@b�2�tk�?
             2@        ������������������������       �                     �?        �       �                    �?ҳ�wY;�?	             1@       �       �                    �?     ��?             0@        ������������������������       �                     @        �       �                 pf&@      �?             $@        ������������������������       �                     @        �       �                  �#@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�Y�R_�?&            �Q@        �       �                    �?ףp=
�?             >@       �       �                    �?ȵHPS!�?             :@       �       �                    �?�S����?             3@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�t����?
             1@       �       �                  ��@8�Z$���?             *@        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                 `fV6@D^��#��?            �D@       �       �                   �A@�q�q�?            �@@       �       �                 ��� @H%u��?             9@        �       �                   �;@և���X�?             @       �       �                   �9@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     2@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                 �?�@PN��T'�?�            �p@        �       �                    �?������?X             b@        �       �                    �?���5��?             �L@       �       �                   �=@      �?             L@       �       �                   �<@:�&���?            �C@       �       �                  ��@$G$n��?            �B@       �       �                   �7@���}<S�?             7@        �       �                   �5@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        
             1@        �       �                 ��(@d}h���?             ,@       �       �                    �?���!pc�?             &@       ������������������������       ��z�G��?             $@        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     1@        ������������������������       �                     �?        �       �                 �{@t��ճC�?8             V@       �       �                   @@@ �Cc}�?$             L@       �       �                    �?�S����?             C@       �       �                    ?@�MI8d�?            �B@       �       �                 ���@(N:!���?            �A@        �       �                 ���@�q�q�?             @       �       �                    �?z�G�z�?             @       �       �                 @33@      �?             @        �       �                    6@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ��@ 	��p�?             =@        ������������������������       �                     *@        �       �                   �4@      �?             0@        ������������������������       �                     &@        �       �                    �?���Q��?             @       �       �                 �1@      �?             @       �       �                   �8@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     2@        ������������������������       �                     @@        �       �                    �?��n��?Y            @_@        �       �                 �yg(@r�q��?             @        �       �                @�µ0@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 @3�@�p�I�?U            �]@        �       �                   �?@�q�q�?             (@        ������������������������       �                     @        �       �                    �?      �?              @       �       �                   �D@և���X�?             @       �       �                   �A@z�G�z�?             @       ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       $                   @pN�Z��?O            �Z@       �                          �?J� ��w�?D             W@       �                       �T)D@�LQ�1	�?2            @Q@       �                          �?     ��?-             P@       �                         �>@@4և���?)             L@       �                          (@dP-���?!            �G@       �                          �:@�����?             E@       �       �                   �3@���7�?             6@        �       �                   �2@ףp=
�?             $@       ������������������������       �                      @        ������������������������       �      �?              @        ������������������������       �        
             (@                                �;@R���Q�?             4@        ������������������������       �                     �?                              ��) @�KM�]�?             3@        ������������������������       �                     "@                              `��!@z�G�z�?             $@        ������������������������       �                     �?                                �<@�����H�?             "@       ������������������������       �                     @        	      
                ���"@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@                              @�$@      �?              @        ������������������������       �                     @                                @7@      �?             @        ������������������������       �                      @        ������������������������       �                      @                                 >@���Q��?             @                                ;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @                                 �?��+7��?             7@                                �?�E��ӭ�?             2@        ������������������������       �                     "@                              `f2@X�<ݚ�?             "@                                �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @               !                   ;@z�G�z�?             @        ������������������������       �                      @        "      #                  @A@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     .@        �t�b� )     h�h*h-K ��h/��R�(KM%KK��h]�BP       `{@      q@     �a@     @e@      =@      @               @      =@       @      <@       @      @              6@       @      6@      �?      @              .@      �?      *@      �?      @      �?      @               @      �?       @               @                      �?      �?             �[@     �d@     �[@     �a@       @     �Z@      �?     �Q@      �?      8@              @      �?      1@      �?      �?              0@             �G@      �?      B@              6@      �?      ,@              @      �?      &@              @      �?      @      �?                      @      [@      B@      :@      @      �?              9@      @       @              7@      @      6@      @      $@              (@      @               @      (@      �?       @              @      �?              �?      @              �?             �T@     �@@               @     �T@      ?@               @     �T@      7@      T@      7@      T@      6@      E@      &@      @      @      @      @              @      @              �?              C@       @      @@       @      2@       @       @       @      �?              �?       @      �?      �?              �?      �?                      �?      0@      @      ,@      @      "@      @      "@      @       @      @      @      @       @      @       @       @       @                       @              �?      �?              @              �?       @               @      �?                      �?      @               @              ,@              @              C@      &@      @              @@      &@      ,@      &@      @      "@      @      @      @       @              �?      @      �?       @      �?       @                      �?       @                      @               @      $@       @       @               @       @       @                       @      2@                      �?       @              �?      7@              3@      �?      @              @      �?             �r@      Z@      Q@      P@      O@      P@      D@      .@      @       @       @       @               @       @      @       @                      @      @             �@@      @      &@              6@      @      2@      @      &@      @              �?      &@      @      &@      @      @              @      @              @      @       @      @                       @              �?      @              @              6@     �H@      @      ;@      @      7@      @      0@      �?      �?              �?      �?               @      .@       @      &@       @                      &@              @              @              @      3@      6@      &@      6@      @      6@      @      @      �?      @      �?                      @       @                      2@       @               @              @             �l@      D@     �`@      *@      I@      @     �H@      @      @@      @      @@      @      5@       @      @       @      @                       @      1@              &@      @       @      @      @      @      �?              @                       @      1@              �?             �T@      @      I@      @      @@      @      ?@      @      ?@      @      @       @      @      �?      @      �?      �?      �?      �?                      �?       @              �?                      �?      ;@       @      *@              ,@       @      &@              @       @      @      �?       @      �?              �?       @              �?                      �?               @      �?              2@              @@             �X@      ;@      �?      @      �?       @               @      �?                      @     @X@      6@      @      @              @      @      @      @      @      @      �?      @      �?      �?                       @      �?              W@      .@     @S@      .@      N@      "@      M@      @      J@      @     �E@      @      C@      @      5@      �?      "@      �?       @              �?      �?      (@              1@      @              �?      1@       @      "@               @       @              �?       @      �?      @               @      �?       @                      �?      @              "@              @       @      @               @       @               @       @               @      @       @      �?              �?       @                       @      1@      @      *@      @      "@              @      @      �?      @      �?                      @      @              @      �?       @               @      �?              �?       @              .@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ��(hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMKhuh*h-K ��h/��R�(KMK��h|�B�R                             !@(����7�?�           @�@               	                   �;@�'N��?#            �N@                                   @�����H�?             B@        ������������������������       �                     *@                                ��*4@�㙢�c�?             7@       ������������������������       �        	             1@                                   @�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        
                           @�q�����?             9@        ������������������������       �                     @                                   �?�����?             3@        ������������������������       �                     "@                                   @���Q��?             $@        ������������������������       �                      @                                ��T?@      �?              @        ������������������������       �                      @        ������������������������       �                     @               �                     @�iz�� �?�           X�@               9                    �?�q�q��?�             r@                                   �?�LQ�1	�?-            @Q@        ������������������������       �                     =@               8                    �?���Q��?             D@              #                  I>@�e����?            �C@                                    �?�8��8��?	             (@        ������������������������       �                      @               "                    �?ףp=
�?             $@              !                   �<@�����H�?             "@                                  �9@�q�q�?             @        ������������������������       �                     �?                                 ���,@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        $       3                    �?X�<ݚ�?             ;@       %       0                    �?D�n�3�?             3@       &       '                    >@�n_Y�K�?	             *@        ������������������������       �                     @        (       )                    A@      �?              @        ������������������������       �                      @        *       -                    �?      �?             @       +       ,                   �I@      �?             @       ������������������������       �                      @        ������������������������       �                      @        .       /                   �E@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        1       2                    6@      �?             @        ������������������������       �                     @        ������������������������       �                     @        4       7                   �C@      �?              @        5       6                 8�P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        :       {                  x#J@&ջ�{��?�            `k@       ;       <                    @H���I�?_            �c@        ������������������������       �                     .@        =       x                    �?��Ok�?X            �a@       >       w                    �?����5�?K            �^@       ?       L                    �?<����l�?I            �]@        @       I                    �?�����?             5@       A       B                 `f�)@�X�<ݺ?             2@        ������������������������       �                     @        C       D                     �?�8��8��?
             (@        ������������������������       �                      @        E       H                    7@ףp=
�?             $@       F       G                    ;@      �?              @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                      @        J       K                   �7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        M       N                   �:@Jm_!'1�?8            �X@        ������������������������       �        
             4@        O       R                   �;@�θ�?.            �S@        P       Q                   �5@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        S       `                   �*@DE��2{�?,            �R@        T       W                 `f�)@�n_Y�K�?             :@        U       V                   @L@�z�G��?             $@       ������������������������       �                     @        ������������������������       �                     @        X       _                    G@     ��?             0@       Y       ^                    C@�q�q�?             (@       Z       [                    =@X�<ݚ�?             "@        ������������������������       �                      @        \       ]                    @@����X�?             @        ������������������������       �                      @        ������������������������       ����Q��?             @        ������������������������       �                     @        ������������������������       �                     @        a       b                 ��$:@�q��/��?            �H@        ������������������������       �        	             0@        c       v                    �?"pc�
�?            �@@       d       u                   �J@     ��?             @@       e       j                 `f�;@�����?             3@        f       g                 03k:@���Q��?             @        ������������������������       �                     �?        h       i                   @B@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        k       l                   @>@d}h���?
             ,@        ������������������������       �                     @        m       n                   �>@�q�q�?             "@        ������������������������       �                      @        o       t                 ��yC@؇���X�?             @       p       q                   �A@      �?             @        ������������������������       �                      @        r       s                   @B@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     *@        ������������������������       �                     �?        ������������������������       �                     @        y       z                    �?���N8�?             5@       ������������������������       �        
             0@        ������������������������       �                     @        |       �                    �?ҐϿ<��?%            �N@       }       ~                 03�a@��p\�?            �D@       ������������������������       �                     <@               �                    �?�θ�?             *@       ������������������������       �                      @        �       �                 ���i@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                 `�iJ@ףp=
�?             4@        ������������������������       �                     �?        �       �                   @@@�}�+r��?             3@        ������������������������       �                     "@        �       �                   @D@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        �       �                    �?��,?S�?�            �v@        �       �                 ��Y7@��
P��?B            @Z@       �       �                    �?�L��7Q�?6            @V@        �       �                   �5@r٣����?            �@@        �       �                 03�@և���X�?             @        ������������������������       �                     �?        �       �                   �2@�q�q�?             @       �       �                 �{&@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?���B���?             :@       �       �                    �?z�G�z�?             9@        �       �                 H�%@����X�?             @        ������������������������       �                      @        �       �                    �?���Q��?             @        ������������������������       �                     �?        �       �                  S�2@      �?             @       �       �                   �<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?r�q��?             2@       �       �                    9@d}h���?             ,@        ������������������������       �                     @        �       �                 �&�@�z�G��?             $@        ������������������������       �                     �?        �       �                 pF @�<ݚ�?             "@       �       �                 �&B@      �?              @       ������������������������       �؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?���>4��?             L@       �       �                   �4@�eP*L��?            �K@        �       �                 @3"@�����H�?             "@       ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �&@
;&����?             G@       �       �                 ��l#@
j*D>�?             :@       �       �                    �?�G��l��?             5@       �       �                   �;@b�2�tk�?
             2@        �       �                   �7@      �?              @       ������������������������       �                     @        �       �                    :@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    I@���Q��?             $@       �       �                 `�X!@؇���X�?             @        ������������������������       �                     @        �       �                  SE"@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �*@��Q��?
             4@        ������������������������       �                     @        �       �                    �?      �?	             ,@       �       �                     @      �?             (@       �       �                 ��Y.@�eP*L��?             &@        ������������������������       �                     @        �       �                 03�1@      �?              @       �       �                    ;@r�q��?             @        �       �                 @3�/@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     0@        �       (                  �<@(L���?�             p@       �       �                    �?Xny��?{            �f@        �       �                    �?������?             >@       �       �                 `v�0@      �?             <@       �       �                    0@r�q��?             8@        ������������������������       �                     �?        �       �                 ��y@�LQ�1	�?             7@        ������������������������       �                     @        �       �                   @@�S����?             3@       �       �                   �7@z�G�z�?             .@        �       �                 ���@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �:@�8��8��?
             (@        ������������������������       �                     �?        �       �                 ���@�C��2(�?	             &@        ������������������������       �                     @        �       �                   @<@r�q��?             @       ������������������������       �z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �2@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ��&@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �                       ��L@�ma�H��?f             c@        �       �                   �8@�J�4�?             I@        �       �                    �?�X�<ݺ?             2@        ������������������������       �                     @        �       �                   �5@��S�ۿ?
             .@        �       �                    4@      �?              @       ������������������������       �                     @        �       �                  s@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �                          �?     ��?             @@                              ��@�+$�jP�?             ;@                                �;@      �?             @        ������������������������       �                      @        ������������������������       �                      @                                 ;@�LQ�1	�?             7@        ������������������������       �                      @              	                   �?z�G�z�?             .@                              03�@      �?              @        ������������������������       �                     �?        ������������������������       �����X�?             @        
                      pf�@؇���X�?             @        ������������������������       �                     @                              �?$@      �?             @       ������������������������       �      �?              @        ������������������������       �                      @                              ��@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @                                 $@X�?٥�?G            �Y@                                 @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                �3@`2U0*��?E             Y@        ������������������������       �                     3@                                �4@H�!b	�?:            @T@                                 �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?                              ���5@p�|�i�?5             S@       ������������������������       �        *            �N@              !                   �?z�G�z�?             .@                                  �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        "      #                   9@"pc�
�?	             &@        ������������������������       �                     @        $      '                   �?      �?              @        %      &                   ;@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     @        )      *                   �?z�G�z�?2            �R@        ������������������������       �                     @        +      0                  �=@��<b���?.            @Q@        ,      /                ���"@      �?              @       -      .                   �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        1      J                   �?��.��?*            �N@       2      I                  @F@���B���?$             J@       3      H                   �?��Sݭg�?            �C@       4      5                �&B@����X�?            �A@        ������������������������       �                     @        6      E                  �D@J�8���?             =@       7      8                   ?@ �o_��?             9@        ������������������������       �                     @        9      B                ��i @�q�q�?             5@       :      A                  �B@      �?	             (@       ;      @                  @@@���Q��?             $@       <      ?                @3�@�q�q�?             @       =      >                P�@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        C      D                �T)D@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        F      G                @3�@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             *@        ������������������������       �                     "@        �t�bh�h*h-K ��h/��R�(KMKKK��h]�B�       �{@      q@      1@      F@      @      @@              *@      @      3@              1@      @       @      @                       @      *@      (@              @      *@      @      "@              @      @       @               @      @       @                      @     pz@     �l@     `b@     �a@      8@     �F@              =@      8@      0@      7@      0@      &@      �?       @              "@      �?       @      �?       @      �?      �?              �?      �?              �?      �?              @              �?              (@      .@      &@       @       @      @      @              @      @               @      @      @       @       @       @                       @      �?      �?              �?      �?              @      @              @      @              �?      @      �?      �?      �?                      �?              @      �?             �^@      X@     �Y@      L@      .@             �U@      L@     �T@      D@     �T@     �B@       @      3@      �?      1@              @      �?      &@               @      �?      "@      �?      @      �?      �?              @               @      �?       @      �?                       @      T@      2@      4@              N@      2@      �?       @      �?                       @     �M@      0@      0@      $@      @      @      @                      @      "@      @      @      @      @      @               @      @       @       @              @       @              @      @             �E@      @      0@              ;@      @      :@      @      *@      @       @      @              �?       @       @      �?              �?       @      &@      @      @              @      @               @      @      �?      @      �?       @              �?      �?              �?      �?              @              *@              �?                      @      @      0@              0@      @              5@      D@      @      C@              <@      @      $@               @      @       @      @                       @      2@       @              �?      2@      �?      "@              "@      �?              �?      "@             @q@     �U@      K@     �I@      C@     �I@       @      9@      @      @      �?               @      @      �?      @              @      �?              �?              @      5@      @      4@       @      @               @       @      @      �?              �?      @      �?       @      �?                       @              �?      @      .@      @      &@              @      @      @      �?               @      @      �?      @      �?      @              �?      �?                      @              �?      >@      :@      >@      9@       @      �?      @               @      �?       @                      �?      6@      8@      .@      &@      $@      &@      @      &@      �?      @              @      �?      @      �?                      @      @      @      @      �?      @               @      �?              �?       @                      @      @              @              @      *@              @      @      @      @      @      @      @      @              @      @      �?      @      �?       @               @      �?                      @       @                      �?      �?      �?      �?                      �?              �?      0@             �k@      B@     @d@      5@      6@       @      5@      @      4@      @              �?      4@      @      @              0@      @      (@      @      �?       @               @      �?              &@      �?      �?              $@      �?      @              @      �?      @      �?      �?              @              �?      @      �?                      @      �?      �?      �?                      �?     �a@      *@      E@       @      1@      �?      @              ,@      �?      @      �?      @              @      �?      @                      �?      @              9@      @      6@      @       @       @               @       @              4@      @       @              (@      @      @       @      �?              @       @      @      �?      @              @      �?      �?      �?       @              @       @      @                       @     �X@      @       @      �?              �?       @              X@      @      3@             @S@      @      @      �?      @                      �?     @R@      @     �N@              (@      @      @      �?      @                      �?      "@       @      @              @       @       @       @              �?       @      �?      @              N@      .@      @              K@      .@      @      @      @       @               @      @                      @     �I@      $@      E@      $@      =@      $@      9@      $@      @              3@      $@      2@      @      @              ,@      @      @      @      @      @       @      @       @       @              �?       @      �?               @      @                       @       @      �?       @                      �?      �?      @              @      �?              @              *@              "@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ���~hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM+huh*h-K ��h/��R�(KM+��h|�B�J                             @�6��l�?�           @�@                                   �?�θ�?            �C@        ������������������������       �                     "@               	                    @�z�G��?             >@                                  @      �?             ,@                               ���W@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        
                           �?      �?             0@                                    @؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?                                   �?�����H�?             "@       ������������������������       �                     @                                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               �                     @b�h�{��?�           �@               %                    �?4�M�f��?�             s@                                   �H@Hn�.P��?N             _@                                 �;@ 5x ��?D            �Z@                                  �7@@4և���?             E@                                   �?���!pc�?             &@        ������������������������       �                     @                                  �'@      �?             @        ������������������������       �                      @                                   �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     ?@        ������������������������       �        +            @P@        !       $                   @I@@�0�!��?
             1@        "       #                 03�3@      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     &@        &       C                 ��D:@T�ue�V�?n            �f@        '       B                    �?$�Z����?0             S@       (       A                 ���+@t�7��?(             O@       )       @                 ��\+@H.�!���?              I@       *       +                     �?     ��?             H@        ������������������������       �                     @        ,       ?                   �*@RB)��.�?            �E@       -       .                    @�θ�?            �C@        ������������������������       �                     @        /       0                   �;@      �?             B@        ������������������������       �        	             ,@        1       8                 `f�)@8�A�0��?             6@       2       7                 `f�&@���!pc�?             &@       3       4                   �H@և���X�?             @       ������������������������       �                     @        5       6                   �P@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        9       >                    G@�eP*L��?             &@       :       ;                   @B@؇���X�?             @        ������������������������       �                     @        <       =                   @D@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     (@        ������������������������       �                     ,@        D       E                 03k:@�#ʆA��?>            �Z@        ������������������������       �                     @        F       c                    �?d,���O�?<            �Y@        G       Z                    �?v�X��?             F@       H       U                   �G@�q�q�?             >@       I       N                    �?��<b���?             7@       J       M                   �;@�t����?             1@        K       L                   �8@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     *@        O       P                 ��3Q@      �?             @        ������������������������       �                     �?        Q       T                   �:@���Q��?             @       R       S                   �5@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        V       Y                    �?����X�?             @       W       X                 ��L@@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        [       `                    �?d}h���?             ,@        \       ]                 h��Q@r�q��?             @        ������������������������       �                     @        ^       _                    6@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        a       b                   @K@      �?              @       ������������������������       �                     @        ������������������������       �                      @        d       e                    �?^l��[B�?'             M@        ������������������������       �                     �?        f       �                   �J@�MWl��?&            �L@       g       �                    �?�^�����?            �E@       h       y                    �?�G�z�?             D@       i       x                     �?      �?             8@       j       q                   �>@�û��|�?             7@        k       p                   @G@�q�q�?             (@       l       o                 `fF<@      �?              @       m       n                   @B@�q�q�?             @        ������������������������       �      �?             @        ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     @        r       w                   �=@�C��2(�?	             &@       s       v                 ��yC@      �?              @        t       u                   �A@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        z       �                 03oY@      �?             0@       {       �                   @K@z�G�z�?
             .@       |       }                   �?@�q�q�?             "@        ������������������������       �                     �?        ~       �                   0F@      �?              @               �                    +@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 `fFJ@�q�q�?             @        ������������������������       �                     �?        �       �                    7@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     ,@        �       "                ��Y7@��*U�?�            �v@       �       �                    �?&��}��?�            �t@        �       �                   �:@p�ݯ��?2             S@        �       �                    �?     ��?             @@       �       �                    �?X�Cc�?             <@        �       �                 �%@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?$��m��?             :@        �       �                  s�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ���@�LQ�1	�?             7@        ������������������������       �                     @        �       �                    �?      �?             4@       �       �                  �#@�t����?             1@       �       �                 pf� @ףp=
�?             $@        �       �                   �9@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �[$@և���X�?             @        ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                     �?        �       �                    9@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�GN�z�?             F@        �       �                 �&B@�nkK�?             7@       �       �                    �?��S�ۿ?
             .@        ������������������������       �                     @        �       �                    �?ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �A@և���X�?             5@       �       �                 `�X!@������?
             .@        �       �                   �;@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        �       �                   �K@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �                          �?����sV�?�            �o@       �                          @@@��V&��?�             k@       �       �                 ��@nS޸��?j             f@        �       �                    �?�eP*L��?             &@        ������������������������       �                     @        �       �                 `f�@����X�?             @       �       �                    6@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                   �>@�/ C-��?d            �d@       �       �                 ��q1@�t����?\             c@       �       �                    �?X�����?Z            �b@        �       �                 H�Z&@R���Q�?             D@       �       �                   �<@�I�w�"�?             C@       �       �                 ���@tk~X��?             B@       �       �                   �7@�d�����?             3@        ������������������������       �                     @        �       �                   �:@      �?	             0@        ������������������������       �                     �?        �       �                 ���@�r����?             .@        ������������������������       �                     @        �       �                   @<@�<ݚ�?             "@       ������������������������       �      �?              @        ������������������������       �                     �?        �       �                    �?�t����?
             1@        ������������������������       �                      @        �       �                  s�@�r����?	             .@        ������������������������       �                     @        �       �                 ��(@"pc�
�?             &@       ������������������������       �z�G�z�?             $@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                   �0@HQ˄�ľ?A            @[@        �       �                 pFD!@և���X�?             @        �       �                 pf�@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 �?$@`'�J�?=            �Y@        �       �                 ��@H%u��?             9@       �       �                    7@���N8�?             5@        ������������������������       �                     &@        �       �                   �8@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        �       �                   �7@      �?             @       ������������������������       �                      @        ������������������������       �                      @        �       �                   �"@�e���@�?-            @S@       ������������������������       �        (            �Q@        �       �                    (@؇���X�?             @        �       �                   �<@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �2@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                 �Y5@�n_Y�K�?             *@        ������������������������       �                     @        �       �                   �?@      �?             $@        ������������������������       �                     �?        �       �                   �@X�<ݚ�?             "@        ������������������������       �                      @        �       �                 �?�@����X�?             @        ������������������������       �                      @        �       �                 ��I @���Q��?             @       ������������������������       ��q�q�?             @        ������������������������       �                      @                              �?�@P���Q�?             D@       ������������������������       �                     :@              
                   �?؇���X�?             ,@                               �B@"pc�
�?
             &@        ������������������������       �                     @              	                @3�@���Q��?             @                               �D@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                 �?�<ݚ�?             B@                                �?��a�n`�?             ?@                                �?      �?             <@                             ��@z�G�z�?             .@        ������������������������       �                     @                              �&�)@      �?              @                             P�@      �?             @                                �9@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                �:@�	j*D�?             *@                                �?և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @              !                  @A@z�G�z�?             @                                 �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        #      *                   �?�}�+r��?             C@        $      %                0�H@r�q��?             (@        ������������������������       �                      @        &      '                   ;@      �?             @        ������������������������       �                     �?        (      )                   >@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     :@        �t�bh�h*h-K ��h/��R�(KM+KK��h]�B�       0{@     Pq@      "@      >@              "@      "@      5@      @      @      �?      @              @      �?              @               @      ,@      �?      @              @      �?              �?       @              @      �?      �?              �?      �?             �z@     �n@     `b@     �c@      @     �]@      @      Z@      @     �C@      @       @              @      @      @               @      @      �?      @                      �?              ?@             @P@      @      ,@      @      @              @      @                      &@     �a@     �D@     @P@      &@     �I@      &@     �C@      &@     �C@      "@      @              A@      "@      >@      "@      @              ;@      "@      ,@              *@      "@       @      @      @      @      @              �?      @              @      �?              @              @      @      �?      @              @      �?       @      �?                       @      @              @                       @      (@              ,@              S@      >@              @      S@      :@      ?@      *@      4@      $@      2@      @      .@       @       @       @       @                       @      *@              @      @              �?      @       @      �?       @      �?                       @       @               @      @       @      @       @                      @              �?      &@      @      @      �?      @               @      �?              �?       @              @       @      @                       @     �F@      *@      �?              F@      *@      >@      *@      ;@      *@      .@      "@      ,@      "@      @       @      @      @      @       @      @      �?      �?      �?               @              @      $@      �?      @      �?       @      �?       @                      �?      @              @              �?              (@      @      (@      @      @      @      �?              @      @      �?      �?              �?      �?              @       @      �?              @       @      @                       @      @                      �?      @              ,@             pq@      V@     `n@     �U@      <@      H@      2@      ,@      2@      $@      �?      �?              �?      �?              1@      "@       @      �?              �?       @              .@       @              @      .@      @      (@      @      "@      �?       @      �?       @                      �?      @              @      @              @      @      �?      �?               @      �?              �?       @              @                      @      $@      A@      �?      6@      �?      ,@              @      �?      "@              "@      �?                       @      "@      (@      @      &@      @      �?              �?      @                      $@      @      �?      @                      �?     �j@      C@     `g@      >@     �b@      <@      @      @      @               @      @       @      @       @                      @               @     �a@      7@     �`@      2@     �`@      0@      ?@      "@      =@      "@      =@      @      ,@      @              @      ,@       @      �?              *@       @      @              @       @      @       @      �?              .@       @       @              *@       @      @              "@       @       @       @      �?                       @       @             �Y@      @      @      @      �?      @      �?                      @      @             �X@      @      6@      @      4@      �?      &@              "@      �?              �?      "@               @       @       @                       @      S@      �?     �Q@              @      �?       @      �?       @                      �?      @               @       @       @                       @       @      @      @              @      @              �?      @      @               @      @       @       @              @       @      �?       @       @              C@       @      :@              (@       @      "@       @      @              @       @      �?       @      �?      �?              �?       @              @              <@       @      8@      @      5@      @      (@      @      @              @      @      �?      @      �?      �?              �?      �?                       @      @              "@      @      @      @              @      @              @              @              @      �?       @      �?              �?       @               @              B@       @      $@       @       @               @       @              �?       @      �?       @                      �?      :@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJCLUhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM9huh*h-K ��h/��R�(KM9��h|�B@N         �                     @Dl���v�?�           @�@                                  �1@d ���T�?�            �s@                                ��f`@ 7���B�?             ;@       ������������������������       �                     9@                                �(\�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               m                  ��T@�d�~V��?�            0r@       	       b                    �?N�R���?�            @n@       
                           @f�Ý��?�            @l@        ������������������������       �                     ,@                                   �?������?�            �j@                                  �H@�}�+r��?,             S@                                  �?��ɉ�?$            @P@       ������������������������       �                    �A@                                   �?��S�ۿ?             >@        ������������������������       �                     "@                                    �?�����?             5@        ������������������������       �                     @                                    @؇���X�?             ,@                                 �7@8�Z$���?             *@        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �                     �?                                �DD@"pc�
�?             &@                                   �?�q�q�?             @                                ���;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @                a                 03�M@� =[y�?W             a@       !       N                    �?��,?S�?N            @^@       "       =                     �?�ZD����?<            @V@       #       $                   �;@     ��?             H@        ������������������������       �                     �?        %       <                    �?p�v>��?            �G@       &       7                   �>@�X����?             F@       '       2                 �ܵ<@*;L]n�?             >@       (       )                   �A@������?             1@        ������������������������       �                     @        *       +                   �E@�q�q�?             (@        ������������������������       �                      @        ,       -                 ��:@z�G�z�?             $@        ������������������������       �                     �?        .       1                    J@�<ݚ�?             "@        /       0                   @G@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        3       4                   �J@�	j*D�?             *@       ������������������������       �                      @        5       6                   @Q@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        8       ;                    �?@4և���?	             ,@        9       :                    G@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     @        >       M                    M@� ��1�?            �D@       ?       @                   �;@8�Z$���?            �C@        ������������������������       �        	             &@        A       B                    �?d}h���?             <@        ������������������������       �                      @        C       D                   �@@8�Z$���?             :@        ������������������������       �                     "@        E       L                    F@������?             1@        F       K                   @C@      �?              @       G       H                   �'@և���X�?             @        ������������������������       �                     �?        I       J                   �3@      �?             @       ������������������������       ����Q��?             @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                      @        O       `                   �C@     ��?             @@       P       _                   �A@��+7��?             7@       Q       X                     �?��s����?             5@        R       S                 `fFJ@      �?              @        ������������������������       �                     @        T       W                 `f�K@      �?             @       U       V                    7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        Y       ^                    :@$�q-�?	             *@       Z       [                   �7@      �?              @       ������������������������       �                     @        \       ]                   �@@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �        	             .@        c       h                   @A@     ��?	             0@       d       g                    �?�C��2(�?             &@        e       f                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        i       l                    @���Q��?             @       j       k                    E@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        n       u                    �?؇���X�?            �H@       o       p                  "�b@@-�_ .�?            �B@       ������������������������       �                     8@        q       t                 Ъ�c@8�Z$���?	             *@        r       s                   �7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        v                        p�w@�q�q�?             (@       w       ~                 �U�^@      �?             $@       x       y                    �?      �?              @        ������������������������       �                     @        z       }                    �?      �?             @       {       |                   �D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?��머��?�            �x@        �       �                    �?6C�z��?G            �\@        �       �                   �"@�q�q�?             E@        ������������������������       �                     @        �       �                    �?p�ݯ��?             C@        �       �                    7@�z�G��?             $@       �       �                 �%@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ��g2@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?      �?             <@       �       �                   �5@���B���?             :@        �       �                  s�@���Q��?             @        ������������������������       �                      @        �       �                 @�@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?؇���X�?             5@       �       �                 ���@r�q��?             2@        ������������������������       �                     �?        �       �                    9@�t����?
             1@        ������������������������       �                     �?        �       �                  s�@      �?	             0@        ������������������������       �                      @        �       �                 �&B@؇���X�?             ,@       ������������������������       �r�q��?             (@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�q�q�?.             R@       �       �                    @�Gi����?            �B@       �       �                    �?<=�,S��?            �A@       �       �                 ���@�P�*�?             ?@        ������������������������       �                     @        �       �                   �>@r�q��?             8@       �       �                   �9@�t����?             1@        �       �                    7@؇���X�?             @       �       �                    5@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 @3�@���Q��?             $@       �       �                 �?�@      �?             @        �       �                   �@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    =@r�q��?             @        ������������������������       �                      @        �       �                 @3#%@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    C@؇���X�?             @        ������������������������       �                     @        �       �                    K@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?4�2%ޑ�?            �A@        �       �                   �@@���Q��?             $@       �       �                   �=@      �?              @       �       �                    ;@�q�q�?             @       �       �                 @3�/@z�G�z�?             @       �       �                   �6@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    @�J�4�?             9@        �       �                 ��T?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �?@�C��2(�?             6@       �       �                    @�}�+r��?             3@       ������������������������       �                     "@        �       �                   �6@ףp=
�?             $@        �       �                 ���3@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   �C@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       0                   �?��W��?�            �q@       �       �                    �?     ��?�             p@        �       �                 �y�#@�חF�P�?             ?@       �       �                    8@ �Cc}�?             <@        �       �                    �?      �?             @       �       �                 �{@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                   @@ �q�q�?             8@       �       �                 ���@��S�ۿ?
             .@        ������������������������       �                     @        �       �                   @<@�����H�?             "@       ������������������������       �r�q��?             @        ������������������������       �                     @        ������������������������       �                     "@        �       �                    7@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                    )@�e�;�?�             l@        ������������������������       �                     @        �       /                   �?���L���?�            @k@       �                         �<@p@T����?r            �g@       �       �                   �4@$�q-�?I            @]@        ������������������������       �                     B@        �                          ;@�����H�?6            @T@        �       �                 @33@r�q��?             >@        ������������������������       �                      @        �                          �9@ �Cc}�?             <@       �       �                 ��L@HP�s��?             9@        �       �                 ���@      �?              @        ������������������������       �                     @        �       �                   �6@      �?             @        �       �                  s@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        
             1@                              d�"@@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?                                @<@�:�]��?!            �I@                             ��) @HP�s��?              I@                                �?���N8�?             E@                               s�@�X�<ݺ?
             2@        ������������������������       �                     @        	      
                ��(@�C��2(�?             &@       ������������������������       �      �?              @        ������������������������       �                     @                               sW@ �q�q�?             8@                              ��@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     4@                              pf� @      �?              @        ������������������������       �                     �?                              �T�C@؇���X�?             @        ������������������������       �                     @        ������������������������       �      �?             @        ������������������������       �                     �?              (                  @@@\�CX�?)            �Q@                                 �?X�<ݚ�?             ;@                                 >@      �?             @        ������������������������       �                     @        ������������������������       �                     �?              '                ���"@
;&����?             7@                               �>@D�n�3�?
             3@        ������������������������       �                     @              "                �?�@�q�q�?             (@               !                  �@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        #      $                  �?@؇���X�?             @        ������������������������       �                     �?        %      &                ��i @r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        )      .                @3�@`���i��?             F@       *      -                  @F@���N8�?             5@        +      ,                   E@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                     7@        ������������������������       �                     >@        1      2                ��A>@ �q�q�?             8@        ������������������������       �                     (@        3      8                   @�8��8��?             (@        4      7                ���A@r�q��?             @        5      6                   @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �t�b��-     h�h*h-K ��h/��R�(KM9KK��h]�B�        {@     `q@      a@     �f@      �?      :@              9@      �?      �?              �?      �?             �`@     �c@      `@     �\@     @_@     @Y@      ,@             �[@     @Y@      @      R@       @     �O@             �A@       @      <@              "@       @      3@              @       @      (@       @      &@       @                      &@              �?       @      "@       @      @       @      �?              �?       @                      @              @     �Z@      =@      W@      =@     �P@      7@     �@@      .@              �?     �@@      ,@      >@      ,@      1@      *@      *@      @      @               @      @               @       @       @      �?              @       @       @       @       @                       @      @              @      "@               @      @      �?      @                      �?      *@      �?       @      �?       @                      �?      &@              @             �@@       @     �@@      @      &@              6@      @               @      6@      @      "@              *@      @      @      @      @      @      �?              @      @       @      @      �?                      �?      "@                       @      :@      @      1@      @      1@      @      @      @      @              �?      @      �?       @      �?                       @              �?      (@      �?      @      �?      @              @      �?              �?      @              @                       @      "@              .@              @      *@      �?      $@      �?      �?              �?      �?                      "@       @      @       @       @       @                       @              �?      @      E@       @     �A@              8@       @      &@       @      �?              �?       @                      $@      @      @      @      @      @      @              @      @      �?      �?      �?              �?      �?               @               @                       @     �r@      X@      L@      M@      ,@      <@              @      ,@      8@      @      @      @      �?              �?      @               @       @       @                       @      @      5@      @      5@       @      @               @       @      �?       @                      �?      @      2@      @      .@      �?               @      .@              �?       @      ,@               @       @      (@       @      $@               @              @       @              E@      >@      .@      6@      *@      6@      *@      2@              @      *@      &@      (@      @      @      �?       @      �?       @                      �?      @              @      @      �?      @      �?      �?              �?      �?                       @      @      �?       @              @      �?      @                      �?      �?      @              @      �?      @      �?                      @              @       @              ;@       @      @      @      @       @      @       @      @      �?      �?      �?      �?                      �?      @                      �?       @                       @      5@      @      �?       @      �?                       @      4@       @      2@      �?      "@              "@      �?       @      �?              �?       @              @               @      �?              �?       @             @n@      C@     `k@     �B@      :@      @      9@      @       @       @      �?       @      �?                       @      �?              7@      �?      ,@      �?      @               @      �?      @      �?      @              "@              �?       @               @      �?              h@      @@              @      h@      9@     `d@      9@      [@      "@      B@              R@      "@      9@      @               @      9@      @      7@       @      @       @      @               @       @      �?      �?      �?                      �?      �?      �?              �?      �?              1@               @      �?       @                      �?     �G@      @      G@      @      D@       @      1@      �?      @              $@      �?      @      �?      @              7@      �?      @      �?      �?               @      �?      4@              @       @              �?      @      �?      @              @      �?      �?             �K@      0@      (@      .@      �?      @              @      �?              &@      (@      &@       @      @              @       @      @       @               @      @              �?      @              �?      �?      @              @      �?                      @     �E@      �?      4@      �?       @      �?       @                      �?      (@              7@              >@              7@      �?      (@              &@      �?      @      �?      �?      �?              �?      �?              @              @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ���hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMUhuh*h-K ��h/��R�(KMU��h|�B@U                              @#�[5]�?�           @�@                                03�;@�!���?             A@                                   �?�X�<ݺ?             2@                                   �?؇���X�?             @                                  �?r�q��?             @        ������������������������       �                      @               
                    �?      �?             @               	                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@                                   @      �?             0@                                �-]@r�q��?             @       ������������������������       �                     @                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   @ףp=
�?             $@                                  @      �?              @        ������������������������       �                     �?                                   �?؇���X�?             @        ������������������������       �                     �?                                   �?r�q��?             @        ������������������������       �                     �?                                ��T?@z�G�z�?             @        ������������������������       �                      @                                   �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        !       &                `fFJ@&�L��?�           0�@       "                        `�X!@@E>���?f           �@        #       2                 ��}@�p ��?�            �n@        $       %                 ��@$Q�q�?(            �O@        ������������������������       �                     5@        &       '                    �?�����?             E@        ������������������������       �                     �?        (       1                    �?��p\�?            �D@       )       *                 ��@�L���?            �B@        ������������������������       �                      @        +       0                    �?��?^�k�?            �A@        ,       -                 ���@P���Q�?             4@       ������������������������       �                     (@        .       /                    8@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     .@        ������������������������       �                     @        3       >                   �3@�s�;�w�?u            �f@        4       5                  s�@b�2�tk�?             2@        ������������������������       �                     @        6       =                     @������?             .@       7       8                 pf�@d}h���?
             ,@        ������������������������       �                     @        9       :                   �0@�z�G��?             $@        ������������������������       ����Q��?             @        ;       <                   �2@z�G�z�?             @       ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     �?        ?       x                   @@@6YE�t�?h            �d@       @       o                   �>@�8����?T            �`@       A       V                    �?��.��?L            �^@        B       U                   �<@�E��ӭ�?             B@       C       L                    �?��R[s�?            �A@        D       E                   �5@�n_Y�K�?	             *@        ������������������������       �                      @        F       G                    9@���!pc�?             &@        ������������������������       �                     �?        H       I                  ��@�z�G��?             $@        ������������������������       �                      @        J       K                 pF @      �?              @       ������������������������       �                     @        ������������������������       �                     �?        M       N                   �8@���7�?             6@        ������������������������       �                     �?        O       P                    �?���N8�?
             5@        ������������������������       �                      @        Q       T                 ��(@$�q-�?             *@       R       S                 03�@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       ������H�?             "@        ������������������������       �                     @        ������������������������       �                     �?        W       j                   �;@X�EQ]N�?7            �U@       X       c                    �?�������?             F@       Y       b                    �?4?,R��?             B@        Z       [                 pf�@      �?              @        ������������������������       �                      @        \       a                   �9@      �?             @       ]       `                 pff@      �?             @       ^       _                   �7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     <@        d       i                    �?      �?              @       e       f                   �6@z�G�z�?             @        ������������������������       �                     �?        g       h                 pff@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        k       l                 ��) @�Ń��̧?             E@       ������������������������       �                    �B@        m       n                 pf� @z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        p       q                 �?�@���|���?             &@        ������������������������       �                      @        r       s                   �?@X�<ݚ�?             "@        ������������������������       �                     �?        t       w                 ��i @      �?              @       u       v                 @3�@և���X�?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     �?        y       z                    �?      �?             @@        ������������������������       �                     @        {       |                 �?�@XB���?             =@       ������������������������       �        	             0@        }       ~                   �E@$�q-�?             *@       ������������������������       �                     (@        ������������������������       �                     �?        �       %                   @���#��?�            �t@       �       �                     @&�bi��?�            �t@       �       �                    �?2��ƾ�?{            @i@       �       �                    �?����T�?w            �h@       �       �                    �?�8 a]��?d            �e@        �       �                   �;@ i���t�?            �H@        �       �                    �?�<ݚ�?	             2@        ������������������������       �                      @        �       �                   �5@      �?             0@        ������������������������       �                     "@        �       �                   �9@և���X�?             @        ������������������������       ����Q��?             @        �       �                   �/@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ���;@�g�y��?             ?@       ������������������������       �                     ;@        �       �                 03�>@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �F@R�f?���?H             _@       �       �                     �?�����?3            �U@        �       �                   �?@X�Cc�?             <@       �       �                    �?���y4F�?             3@        ������������������������       �                     @        �       �                    �?      �?	             0@       �       �                 `f�D@����X�?             ,@       �       �                   �;@���Q��?             $@        ������������������������       �                     �?        �       �                   �<@�q�q�?             "@       �       �                   �A@և���X�?             @       �       �                   `@@z�G�z�?             @       �       �                 `f�<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                 `f�<@�q�q�?             "@       ������������������������       �      �?             @        ������������������������       �                     @        �       �                   @D@�^����?%            �M@       �       �                   �*@4��?�?!             J@       �       �                 `fF)@      �?             @@        �       �                   �5@@4և���?	             ,@        �       �                    &@؇���X�?             @       �       �                   �1@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �      �?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �;@r�q��?             2@        ������������������������       �                     @        �       �                    =@���!pc�?             &@        ������������������������       �                     �?        �       �                    @@z�G�z�?             $@        ������������������������       �                     @        �       �                   @B@�q�q�?             @       ������������������������       ��q�q�?             @        ������������������������       �                     @        �       �                    �?P���Q�?             4@        ������������������������       �                     @        �       �                   �@@@4և���?	             ,@        �       �                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        �       �                   �3@����X�?             @        ������������������������       ��q�q�?             @        ������������������������       �                     @        �       �                   �N@@-�_ .�?            �B@       �       �                    �?      �?             @@       �       �                   �H@XB���?             =@        �       �                     �?ףp=
�?             $@       �       �                   �G@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        
             3@        ������������������������       �                     @        �       �                 `f�2@z�G�z�?             @        �       �                   �P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?r�q��?             8@        ������������������������       �        	             (@        �       �                   pA@�8��8��?
             (@       ������������������������       �                      @        �       �                    �?      �?             @        ������������������������       �                     �?        �       �                   �B@�q�q�?             @       �       �                    +@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �                          �?0,Tg��?K            �_@       �                          �?�x�(��?:             W@        �       �                    7@�eP*L��?             F@        �       �                    �?���!pc�?             &@       �       �                    �?�z�G��?             $@       �       �                    �?r�q��?             @        ������������������������       �                      @        �       �                  �#@      �?             @        ������������������������       �                      @        �       �                 �[$@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ��'@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        �                           �?���|���?            �@@        �       �                   �;@d}h���?             ,@        ������������������������       �                     @        �       �                  SE"@�z�G��?             $@        ������������������������       �                     @        �       �                  S�2@և���X�?             @       �       �                  S�(@      �?             @        �       �                    I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �<@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?                              03�1@�\��N��?             3@                                �?z�G�z�?             $@                             ���(@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?              
                   �?�<ݚ�?             "@             	                   �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @                                 �?8��8���?             H@                                 ;@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                 �?�����H�?            �F@        ������������������������       �                     $@                                 ,@؇���X�?            �A@        ������������������������       �                     @                              ���#@�g�y��?             ?@                                �<@ףp=
�?             $@       ������������������������       �                      @                                 C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     5@              $                03�7@�IєX�?             A@                                 7@"pc�
�?             &@        ������������������������       �                     @                                 �?      �?              @        ������������������������       �                     �?               #                  @A@؇���X�?             @       !      "                   �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     7@        ������������������������       �                     @        '      T                   @�JY�8��?@             Y@       (      K                   �?Bԅ���?<            �W@       )      0                   �?2X��ʑ�?5            �U@       *      +                ���a@`'�J�?            �I@       ������������������������       �                    �A@        ,      /                03c@      �?             0@        -      .                   �?�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     $@        1      J                  �B@����X�?            �A@       2      9                   �?X�Cc�?             <@        3      8                �̾w@�q�q�?             (@       4      5                  �8@�����H�?             "@        ������������������������       �                     @        6      7                   :@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        :      I                03�X@      �?
             0@       ;      @                   �?����X�?	             ,@        <      ?                ��P@�q�q�?             @       =      >                   >@���Q��?             @       ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                     �?        A      H                  �@@      �?              @       B      G                   >@���Q��?             @       C      F                   <@      �?             @       D      E                   7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        L      S                    �?X�<ݚ�?             "@       M      N                   �?�q�q�?             @        ������������������������       �                     @        O      P                ���[@�q�q�?             @        ������������������������       �                     �?        Q      R                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �t�bh�h*h-K ��h/��R�(KMUKK��h]�BP       �}@     �m@      &@      7@      �?      1@      �?      @      �?      @               @      �?      @      �?      �?      �?                      �?               @              �?              &@      $@      @      �?      @              @      �?      �?      �?                      �?      "@      �?      @      �?      �?              @      �?      �?              @      �?      �?              @      �?       @               @      �?       @                      �?       @             }@     �j@     �z@     �b@     @j@      B@     �M@      @      5@              C@      @              �?      C@      @      A@      @               @      A@      �?      3@      �?      (@              @      �?              �?      @              .@              @             �b@      @@      &@      @              @      &@      @      &@      @      @              @      @      @       @      @      �?      @              �?      �?              �?     �a@      9@     @[@      8@     �Y@      4@      :@      $@      :@      "@      @       @       @              @       @              �?      @      @       @              �?      @              @      �?              5@      �?      �?              4@      �?       @              (@      �?      "@      �?      �?               @      �?      @                      �?      S@      $@     �A@      "@      ?@      @      @      @               @      @      @      @      �?      �?      �?              �?      �?               @                       @      <@              @      @      �?      @              �?      �?      @              @      �?              @             �D@      �?     �B@              @      �?              �?      @              @      @       @              @      @              �?      @      @      @      @      @       @              �?      �?              ?@      �?      @              <@      �?      0@              (@      �?      (@                      �?     @k@     �\@     �j@     �\@     @^@     @T@     @^@      S@     �[@     �O@      @      F@      @      ,@               @      @      (@              "@      @      @      @       @      �?      �?              �?      �?              �?      >@              ;@      �?      @      �?                      @     @Z@      3@     �Q@      1@      2@      $@      .@      @      @              (@      @      $@      @      @      @              �?      @      @      @      @      @      �?      �?      �?      �?                      �?      @                       @       @              @               @              @      @      @      �?              @      J@      @     �G@      @      <@      @      *@      �?      @      �?      @      �?      �?              @      �?       @              @              .@      @      @               @      @              �?       @       @      @              @       @      �?       @      @              3@      �?      @              *@      �?      @      �?      @                      �?      "@              @       @      �?       @      @             �A@       @      ?@      �?      <@      �?      "@      �?      @      �?      @                      �?       @              3@              @              @      �?      �?      �?              �?      �?              @              &@      *@              (@      &@      �?       @              @      �?      �?               @      �?      �?      �?              �?      �?              �?                      @     @W@     �@@     �N@      ?@      4@      8@       @      @      @      @      @      �?       @              @      �?       @              �?      �?              �?      �?               @       @               @       @              �?              (@      5@      @      &@              @      @      @              @      @      @      @      @      �?      �?      �?                      �?       @       @       @                       @              �?      "@      $@       @       @      �?       @      �?                       @      �?              @       @      @       @      @                       @      @             �D@      @      �?       @               @      �?              D@      @      $@              >@      @              @      >@      �?      "@      �?       @              �?      �?              �?      �?              5@              @@       @      "@       @      @              @       @              �?      @      �?      @      �?      @                      �?      @              7@              @             �B@     �O@      @@     �O@      ;@     �M@       @     �H@             �A@       @      ,@       @      @              @       @                      $@      9@      $@      2@      $@       @      @       @      �?      @              @      �?              �?      @                      @      $@      @      $@      @      @       @      @       @      @      �?              �?      �?              @       @      @       @      @      �?      �?      �?      �?                      �?       @                      �?      @                       @      @              @      @       @      @              @       @      �?      �?              �?      �?              �?      �?              @              @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ"�a,hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM)huh*h-K ��h/��R�(KM)��h|�B@J                             @�6��l�?�           @�@                                   �?�^�����?            �E@        ������������������������       �                     "@                                   @h+�v:�?             A@                               �-]@��2(&�?             6@                                 �&@�}�+r��?             3@        ������������������������       �                     �?        ������������������������       �                     2@        	       
                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                   �?r�q��?             (@        ������������������������       �                     @                                   @�q�q�?             @                               ��T?@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?               (                   @`S�as��?�           �@              �                    �? n1U�5�?�           8�@              ^                    �?�!�a�?,           p|@               !                    �?z�G�z�?[            �`@                                 hލC@8�Z$���?             :@                                `v7<@���|���?	             &@                                   @�<ݚ�?             "@        ������������������������       �                      @                                H�%@����X�?             @        ������������������������       �                     @                                   �?      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        	             .@        "       U                   �=@:䠍[O�?I            @[@       #       ,                     @�(�Tw��?2            �S@        $       %                    �? 7���B�?             ;@        ������������������������       �                     �?        &       +                    �? ��WV�?             :@       '       *                   �3@�IєX�?
             1@        (       )                   �9@�����H�?             "@        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@        -       J                 @3�@j���� �?!            �I@       .       /                    @����>�?            �B@        ������������������������       �                     �?        0       I                    �?      �?             B@       1       :                    �?H�V�e��?             A@        2       3                 ���@؇���X�?
             ,@        ������������������������       �                     �?        4       9                 �&B@$�q-�?	             *@       5       6                    9@�����H�?             "@        ������������������������       �                     �?        7       8                 ���@      �?              @        ������������������������       �                      @        ������������������������       �r�q��?             @        ������������������������       �                     @        ;       <                    0@      �?             4@        ������������������������       �                     �?        =       @                   �3@���y4F�?
             3@        >       ?                 P��@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        A       B                   �6@؇���X�?             ,@        ������������������������       �                     @        C       H                   �9@����X�?             @       D       G                    8@�q�q�?             @       E       F                 @3�@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        K       R                    �?d}h���?
             ,@       L       M                    �?�C��2(�?             &@        ������������������������       �                     �?        N       O                  �#@ףp=
�?             $@       ������������������������       �                      @        P       Q                 �[$@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        S       T                 @3�2@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        V       ]                    �?�g�y��?             ?@       W       X                   @B@���7�?             6@       ������������������������       �        	             *@        Y       Z                     @�����H�?             "@       ������������������������       �                     @        [       \                    I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        _       �                    �?أp=
��?�             t@       `       y                     �?����ak�?�            �s@        a       x                 p�w@^(��I�?$            �K@       b       k                    �?�T`�[k�?#            �J@        c       j                 `f�B@R���Q�?             4@       d       e                 ���<@�z�G��?             $@        ������������������������       �                     @        f       i                 ��>@      �?             @        g       h                   �E@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        l       m                 `fF:@���!pc�?            �@@        ������������������������       �                     @        n       u                   �J@$��m��?             :@       o       t                   �>@X�<ݚ�?             2@       p       s                   @>@�q�q�?             (@       q       r                   �B@���Q��?             $@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        v       w                    R@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        z       �                 0��D@��0���?�            p@       {       �                    �?`0�Ƒg�?�            �o@        |       }                   �7@�<ݚ�?             B@        ������������������������       �                     @        ~       �                 83�0@6YE�t�?            �@@              �                 ���@      �?             @@        ������������������������       �                     &@        �       �                 �R,@��s����?             5@       �       �                     @�<ݚ�?             2@        ������������������������       �                     �?        �       �                   �<@@�0�!��?
             1@       �       �                   @<@؇���X�?             ,@       �       �                   @@r�q��?             (@       ������������������������       �"pc�
�?             &@        ������������������������       �                     �?        ������������������������       �                      @        �       �                    ?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                 ��y @ċ��s�?�             k@       �       �                    �?ȵHPS!�?c            �c@        ������������������������       �                     2@        �       �                    1@�LQ�1	�?X            @a@        �       �                 pf�@և���X�?             @        ������������������������       �                      @        ������������������������       �z�G�z�?             @        �       �                 ��) @A5Xo�?U            ``@       �       �                   �>@ףp=
�?T            @`@       �       �                     @`��F:u�?;            �U@        ������������������������       �                     @        �       �                   �;@������?8            �T@       �       �                   �:@HP�s��?"             I@       �       �                 �?$@ �q�q�?              H@        ������������������������       �        	             &@        �       �                 �1@@-�_ .�?            �B@        �       �                   �5@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �3@      �?             @@        �       �                 �?�@      �?             @        ������������������������       �                      @        ������������������������       �      �?              @        ������������������������       �                     <@        ������������������������       �                      @        ������������������������       �                     @@        �       �                   @@@RB)��.�?            �E@        �       �                   �?@      �?             ,@        �       �                 pff@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �@      �?             $@        ������������������������       �                     @        �       �                 @3�@����X�?             @       �       �                 �?�@r�q��?             @        ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                     �?        �       �                   @C@ 	��p�?             =@        ������������������������       �                     .@        �       �                 P�@؇���X�?
             ,@        ������������������������       �                     @        �       �                   �G@�<ݚ�?             "@        �       �                   �D@���Q��?             @       ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                     @��v$���?*            �N@        ������������������������       �                     >@        �       �                 ���"@�g�y��?             ?@        ������������������������       �        
             2@        �       �                    (@$�q-�?             *@        �       �                   �<@z�G�z�?             @       ������������������������       �                     @        �       �                    ?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                     @      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                      @        �       �                    �?      �?y             h@       �       �                 м�9@r٣����?B            �X@        �       �                     @��Zy�?            �C@        ������������������������       �                      @        �       �                    @`՟�G��?             ?@       �       �                    �?��
ц��?             :@        �       �                    �?z�G�z�?             $@       �       �                   @5@�q�q�?             @        ������������������������       �                     �?        �       �                    �?z�G�z�?             @       �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?      �?             0@       �       �                   �6@      �?             $@        ������������������������       �                      @        �       �                 03�1@      �?              @       �       �                   �D@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?r�q��?             @       �       �                   �>@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�?�P�a�?'             N@       �       �                   �8@$�q-�?              J@        ������������������������       �        	             0@        �       �                    ;@�����H�?             B@        �       �                 ���V@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ��H@�FVQ&�?            �@@        �       �                   �E@"pc�
�?             &@       �       �                    @ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     6@        �       �                     @      �?              @       ������������������������       �                     @        ������������������������       �                     @        �                        x#J@��a�n`�?7            @W@       �       �                    �?�C��2(�?(            �P@        ������������������������       �                     (@        �                           )@�����H�?!             K@        ������������������������       �                     @                                �8@�IєX�?            �I@        ������������������������       �                     2@                                �9@�C��2(�?            �@@                                  @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                 �?(;L]n�?             >@             	                м�6@���N8�?             5@       ������������������������       �        	             ,@        
                          �?؇���X�?             @        ������������������������       �                     @                                �:@      �?             @                               �@@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@                                 �?X�<ݚ�?             ;@                             0�"K@     ��?	             0@        ������������������������       �                     �?                                 �?������?             .@                             ���S@�z�G��?             $@        ������������������������       �                     @                                @C@���Q��?             @        ������������������������       �                      @                              @�pX@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                              ��<R@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @               !                   �?���|���?             &@        ������������������������       �                     �?        "      '                   @���Q��?             $@       #      &                    @X�<ݚ�?             "@       $      %                  @F@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     6@        �t�bh�h*h-K ��h/��R�(KM)KK��h]�B�       0{@     Pq@      *@      >@              "@      *@      5@      @      3@      �?      2@      �?                      2@       @      �?       @                      �?      $@       @      @              @       @      @       @      @                       @      �?             `z@     �n@      y@     �n@      s@     �b@      ;@      [@      @      6@      @      @       @      @               @       @      @              @       @       @       @                       @       @                      .@      7@     �U@      6@      L@      �?      :@              �?      �?      9@      �?      0@      �?       @      �?      �?              @               @              "@      5@      >@      $@      ;@      �?              "@      ;@      @      ;@       @      (@      �?              �?      (@      �?       @              �?      �?      @               @      �?      @              @      @      .@      �?              @      .@       @      @              @       @               @      (@              @       @      @       @      �?      �?      �?              �?      �?              �?                      @       @              &@      @      $@      �?      �?              "@      �?       @              �?      �?              �?      �?              �?       @               @      �?              �?      >@      �?      5@              *@      �?       @              @      �?      �?      �?                      �?              "@     Pq@     �E@     �p@     �E@     �D@      ,@     �D@      (@      1@      @      @      @      @              �?      @      �?      �?              �?      �?                       @      $@              8@      "@      @              1@      "@      $@       @      @       @      @      @      @                      @               @      @              @      �?      @                      �?               @     �l@      =@     @l@      ;@      <@       @              @      <@      @      <@      @      &@              1@      @      ,@      @              �?      ,@      @      (@       @      $@       @      "@       @      �?               @               @      �?              �?       @              @                      �?     �h@      3@     @a@      2@      2@              ^@      2@      @      @       @              �?      @     @]@      ,@     @]@      *@     �T@      @      @             �S@      @      G@      @      G@       @      &@             �A@       @      @      �?              �?      @              ?@      �?      @      �?       @              �?      �?      <@                       @      @@              A@      "@      @      @       @       @       @                       @      @      @              @      @       @      @      �?      @               @      �?              �?      ;@       @      .@              (@       @      @              @       @      @       @      @      �?              �?      @                      �?      N@      �?      >@              >@      �?      2@              (@      �?      @      �?      @              �?      �?              �?      �?               @               @       @      �?              �?       @       @              X@      X@      8@     �R@      1@      6@               @      1@      ,@      (@      ,@       @       @       @      @      �?              �?      @      �?       @      �?                       @               @              @      $@      @      @      @       @              @      @      �?      @              @      �?               @              @      �?      @      �?      @                      �?      �?              @              @     �J@      @      H@              0@      @      @@       @      �?              �?       @               @      ?@       @      "@      �?      "@              "@      �?              �?                      6@      @      @              @      @              R@      5@      N@      @      (@              H@      @              @      H@      @      2@              >@      @      �?       @      �?                       @      =@      �?      4@      �?      ,@              @      �?      @              @      �?       @      �?              �?       @              �?              "@              (@      .@      @      &@      �?              @      &@      @      @              @      @       @       @              �?       @               @      �?              �?      @      �?                      @      @      @      �?              @      @      @      @      @      @              @      @               @              �?              6@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�8�hhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM=huh*h-K ��h/��R�(KM=��h|�B@O         �                     @���x�W�?�           @�@               [                  x#J@te��e��?�            �s@              N                    �?�ҹ��?�            �i@                                  @�&!��?k            �e@        ������������������������       �                     *@               M                 �D�H@d ���T�?d            �c@                                  �?��&T)��?_            �b@               	                    4@X�<ݚ�?             ;@        ������������������������       �                      @        
                           �?�q�����?             9@        ������������������������       �                      @                                   =@�t����?             1@                                 �<@�C��2(�?             &@                                   �?؇���X�?             @        ������������������������       �                      @                                  �9@z�G�z�?             @        ������������������������       �                      @                                ���,@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                   A@�q�q�?             @        ������������������������       �                     @                                  �B@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                   �?�g;aS�?N             _@        ������������������������       �                    �A@               4                     �?��f��?:            @V@               1                    K@��}*_��?             ;@              0                   �G@�\��N��?             3@               !                 ��$:@j���� �?             1@        ������������������������       �                      @        "       +                   �E@��S���?             .@       #       $                 03k:@���Q��?             $@        ������������������������       �                     @        %       *                   �A@և���X�?             @       &       '                   @>@z�G�z�?             @        ������������������������       �                      @        (       )                   �>@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ,       /                   �F@z�G�z�?             @       -       .                 `f?@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        2       3                 `fF<@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        5       J                   @N@��� ��?$             O@       6       C                    �?�j��b�?"            �M@       7       B                   �*@HP�s��?             I@       8       =                 `f�)@��-�=��?            �C@        9       <                   �6@��S�ۿ?
             .@        :       ;                   �2@z�G�z�?             @        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     $@        >       ?                   �=@      �?             8@       ������������������������       �                     ,@        @       A                   @B@�z�G��?             $@        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     &@        D       E                   �7@�<ݚ�?             "@        ������������������������       �                     @        F       I                   �B@���Q��?             @        G       H                   �<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        K       L                   �P@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        O       P                    �?     ��?             @@       ������������������������       �                     3@        Q       R                   `6@�	j*D�?             *@        ������������������������       �                      @        S       V                    :@"pc�
�?	             &@        T       U                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        W       Z                    �?�����H�?             "@        X       Y                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        \       �                    �?�ψX�F�?C            @\@       ]       r                 03?U@8�B�q�?8            �W@       ^       a                   �;@Fx$(�?             I@        _       `                    �?$�q-�?	             *@       ������������������������       �                     (@        ������������������������       �                     �?        b       c                    �?��+��?            �B@        ������������������������       �        	             (@        d       e                 �K@ �o_��?             9@        ������������������������       �                      @        f       q                   �L@��<b���?             7@       g       p                     �?؇���X�?             5@       h       i                    �?R���Q�?
             4@        ������������������������       �                     @        j       k                   �G@�θ�?             *@       ������������������������       �                     @        l       m                 p"�P@      �?             @        ������������������������       �                      @        n       o                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        s       |                    �?���V��?            �F@       t       {                    �?�8��8��?             B@       u       z                    �?�S����?             3@       v       w                 ��`g@�IєX�?
             1@       ������������������������       �                     *@        x       y                   �?@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     1@        }       ~                   �?@X�<ݚ�?             "@        ������������������������       �                      @               �                    �?����X�?             @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    4@�X�<ݺ?             2@        �       �                    2@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     *@        �       �                    �?Ҍ�����?�            �x@        �       �                    �?X�<ݚ�?L            @]@       �       �                    �?fK!���?;            �V@       �       �                    �?B�
k���?/            �P@        �       �                 03�@ �o_��?             9@        ������������������������       �                     @        �       �                    �?"pc�
�?             6@        �       �                 H�%@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                 ���@��S�ۿ?             .@        ������������������������       �                     �?        ������������������������       �                     ,@        �       �                     @�D����?             E@       �       �                    �?�99lMt�?            �C@       �       �                    K@���@M^�?             ?@       �       �                 ���@d��0u��?             >@        ������������������������       �                     @        �       �                 ��&@l��
I��?             ;@       �       �                 �[$@R�}e�.�?             :@       �       �                   �;@�X����?             6@       �       �                  �#@���Q��?
             .@       �       �                   �9@�	j*D�?	             *@       �       �                    5@ףp=
�?             $@        ������������������������       �                     @        �       �                  � @      �?             @        �       �                   �7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                   �>@؇���X�?             @       ������������������������       �                     @        �       �                    C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ��Y.@      �?              @        ������������������������       �                     @        �       �                   �=@���Q��?             @       �       �                    9@�q�q�?             @        ������������������������       �                     �?        �       �                    ;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    @      �?             8@       �       �                    �?���Q��?
             4@        �       �                 83�0@      �?              @        ������������������������       �                     @        ������������������������       �                     @        �       �                 P��%@�q�q�?             (@        ������������������������       �                     @        �       �                 `fV6@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    A@���B���?             :@       �       �                   �<@      �?             4@       �       �                    @@�0�!��?             1@       �       �                    @      �?
             0@        �       �                 ��T?@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �                     �?        �       �                    @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �                          �?�7��ެ�?�            `q@       �                       ��q1@�r����?�            @j@       �       �                   �0@,�8����?�            `i@        ������������������������       �                     @        �       �                 �Y�@ףp=
�?�             i@        �       �                   �8@�<ݚ�?             B@        �       �                    5@���|���?             &@       �       �                   �3@�q�q�?             @        ������������������������       �                     �?        �       �                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                 ���@`2U0*��?             9@       ������������������������       �                     5@        �       �                   @<@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        �                          �?��p\�?k            �d@       �       �                   �<@��(\���?h             d@       �       �                    �?������?E             [@        ������������������������       �        
             0@        �       �                    ;@hl �&�?;             W@       �       �                 @3�@ �Jj�G�?"            �K@        ������������������������       �                     =@        �       �                 ��Y @ ��WV�?             :@        �       �                    4@      �?              @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     2@        �       �                   @<@@-�_ .�?            �B@       �       �                 �?$@�X�<ݺ?             B@        �       �                 ��@z�G�z�?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        �       �                 ��) @�g�y��?             ?@       ������������������������       �                     7@        �       �                 pf� @      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �                          �?D>�Q�?#             J@        �                          �?z�G�z�?             .@        �                       �� @؇���X�?             @       �                           ?@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @                                 >@      �?              @        ������������������������       �                      @        ������������������������       �                     @                              @3�@�MI8d�?            �B@                               �C@���N8�?             5@                               �B@�t����?             1@       	      
                �&B@d}h���?
             ,@        ������������������������       �                     @                                @@@�z�G��?             $@                               �@      �?             @        ������������������������       �                      @                              �?�@      �?             @        ������������������������       �                      @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                     @                                �=@      �?             0@                              �̌!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             ,@        ������������������������       �                     @                                 ;@����X�?             @        ������������������������       �                     @                                 >@      �?             @       ������������������������       �                      @        ������������������������       �                      @              2                ��Y7@�������?(             Q@              '                   �?F�����?            �F@        !      "                   7@���!pc�?             &@        ������������������������       �                     @        #      $                   �?      �?             @        ������������������������       �                      @        %      &                 �v6@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        (      1                   �?�������?             A@       )      *                   *@��X��?             <@        ������������������������       �                     @        +      ,                   3@�����?             5@        ������������������������       �                     "@        -      0                pf�'@r�q��?	             (@        .      /                ��@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        3      4                   �?�nkK�?             7@        ������������������������       �                     &@        5      <                   @�8��8��?             (@       6      ;                   @      �?              @       7      8                ��T?@r�q��?             @        ������������������������       �                     @        9      :                   @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �t�b� .     h�h*h-K ��h/��R�(KM=KK��h]�B�       P{@     0q@     �a@      f@     @\@     �V@      Z@      Q@      *@             �V@      Q@     �T@      Q@      (@      .@               @      (@      *@               @      (@      @      $@      �?      @      �?       @              @      �?       @               @      �?              �?       @              @               @      @              @       @      �?              �?       @             �Q@     �J@             �A@     �Q@      2@      1@      $@      $@      "@      $@      @       @               @      @      @      @              @      @      @      @      �?       @               @      �?              �?       @                       @      @      �?       @      �?      �?      �?      �?               @                       @      @      �?      @                      �?      K@       @     �J@      @      G@      @     �A@      @      ,@      �?      @      �?      @              �?      �?      $@              5@      @      ,@              @      @      �?      @      @              &@              @       @      @              @       @      �?       @      �?                       @       @              �?       @               @      �?               @              "@      7@              3@      "@      @               @      "@       @      �?      �?      �?                      �?       @      �?       @      �?              �?       @              @              ;@     �U@      :@     @Q@      3@      ?@      �?      (@              (@      �?              2@      3@              (@      2@      @               @      2@      @      2@      @      1@      @      @              $@      @      @              @      @       @              �?      @              @      �?              �?                       @      @      C@      @     �@@      @      0@      �?      0@              *@      �?      @      �?                      @       @                      1@      @      @       @               @      @       @      �?              �?       @                      @      �?      1@      �?      @              @      �?                      *@     �r@     �X@     @P@      J@      F@     �G@      @@     �A@      @      2@      @              @      2@      @      @              @      @              �?      ,@      �?                      ,@      9@      1@      9@      ,@      3@      (@      3@      &@              @      3@       @      3@      @      .@      @      "@      @      "@      @      "@      �?      @              @      �?      �?      �?              �?      �?               @                      @               @      @      �?      @              �?      �?              �?      �?              @                      �?              �?      @       @      @              @       @      �?       @              �?      �?      �?      �?                      �?       @                      @      (@      (@       @      (@      @      @      @                      @      @      @      @               @      @              @       @              @              5@      @      .@      @      ,@      @      ,@       @      @       @      @                       @      $@                      �?      �?       @               @      �?              @              m@      G@     �f@      <@     �f@      7@              @     �f@      4@      <@       @      @      @      @       @      �?              @       @               @      @                      @      8@      �?      5@              @      �?       @      �?      �?              c@      (@     �b@      (@     @Z@      @      0@             @V@      @      K@      �?      =@              9@      �?      @      �?      �?      �?      @              2@             �A@       @      A@       @      @      �?       @               @      �?      >@      �?      7@              @      �?              �?      @              �?             �E@      "@      (@      @      @      �?      @      �?              �?      @               @              @       @               @      @              ?@      @      0@      @      (@      @      &@      @      @              @      @      @      @               @      @      �?       @              �?      �?      @              �?       @      @              .@      �?      �?      �?      �?                      �?      ,@              @               @      @              @       @       @       @                       @      I@      2@      <@      1@      @       @              @      @      @       @              �?      @      �?                      @      9@      "@      3@      "@              @      3@       @      "@              $@       @       @       @       @                       @       @              @              6@      �?      &@              &@      �?      @      �?      @      �?      @              �?      �?              �?      �?               @              @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJP�dhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM3huh*h-K ��h/��R�(KM3��h|�B�L         d                    �?~�Я��?�           @�@               _                    @��mo*�?�            �m@              .                   �:@��z����?�            �k@               	                    �?<)�%�w�?7            @W@                                033.@8�Z$���?             :@                                pFt*@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        
             3@        
       )                    �?�Z4���?(            �P@              (                 �̌3@��N`.�?!            �K@              #                   �8@��
ц��?            �C@                                  3@����"�?             =@                                   1@r�q��?             @        ������������������������       �                      @                                �y� @      �?             @        ������������������������       �                     �?        ������������������������       �                     @               "                    �?\X��t�?             7@                               ���@�ՙ/�?             5@        ������������������������       �                     @                                ��Y#@��.k���?
             1@                               pff@���Q��?             $@                                   �?�q�q�?             @                                 �5@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @               !                     @����X�?             @                                  �'@r�q��?             @        ������������������������       �                      @        ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                      @        $       '                    �?�z�G��?             $@       %       &                 �&B@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     0@        *       +                     @�q�q�?             (@        ������������������������       �                     @        ,       -                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     @        /       H                    �?      �?S             `@       0       G                    @�L���?1            �R@       1       2                     @�X�<ݺ?/             R@       ������������������������       �                     �I@        3       >                    �?��s����?             5@       4       ;                   �B@�r����?
             .@       5       6                    �?�C��2(�?             &@       ������������������������       �                     @        7       8                 @3�@      �?             @        ������������������������       �                      @        9       :                    =@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        <       =                 `fV!@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ?       @                 ��"@�q�q�?             @        ������������������������       �                     �?        A       F                    �?z�G�z�?             @       B       E                  S�2@�q�q�?             @       C       D                   �<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        I       P                    �?�+$�jP�?"             K@        J       O                   �>@�X�<ݺ?             2@        K       L                     @�����H�?             "@        ������������������������       �                     @        M       N                 pF�-@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        Q       X                    @@      �?             B@        R       S                   �<@      �?             $@        ������������������������       �                     @        T       W                    �?r�q��?             @        U       V                    6@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        Y       Z                   �B@8�Z$���?             :@        ������������������������       �                      @        [       ^                    @�<ݚ�?             2@       \       ]                     @��S�ۿ?
             .@       ������������������������       �        	             ,@        ������������������������       �                     �?        ������������������������       �                     @        `       a                      @������?             .@        ������������������������       �                      @        b       c                   �>@8�Z$���?	             *@       ������������������������       �                     &@        ������������������������       �                      @        e       �                     �?ꀕ<u�?%           �}@        f       }                   �>@D�]�+��?7            �X@        g       |                   �J@X�<ݚ�?            �F@       h       q                    ?@4�B��?            �B@        i       p                   �<@"pc�
�?             &@       j       m                    �?�<ݚ�?             "@        k       l                 �ܵ<@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        n       o                 `f�<@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        r       {                   �G@ȵHPS!�?             :@       s       t                    �?@�0�!��?             1@        ������������������������       �                     @        u       z                    G@�θ�?             *@       v       y                   @D@�C��2(�?             &@        w       x                 ��I*@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                      @        ~       �                    >@r�z-��?"            �J@               �                   �9@�q�q�?             8@        ������������������������       �                     @        �       �                    �?      �?
             4@        �       �                   �;@r�q��?             @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �A@����X�?             ,@        ������������������������       �                     @        �       �                   �<@      �?              @       �       �                   �;@z�G�z�?             @        ������������������������       �                     �?        �       �                   �E@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?П[;U��?             =@        �       �                   @D@�q�q�?             "@        ������������������������       �                     @        �       �                  �}S@      �?             @        ������������������������       �                      @        �       �                    �?      �?             @        ������������������������       �                     �?        �       �                 `��W@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    D@��Q��?             4@        �       �                   @B@�q�q�?             @       �       �                    �?      �?             @       �       �                   �@@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ���[@d}h���?
             ,@       ������������������������       �                     "@        �       �                 `f�h@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                 �?�@4z�_�\�?�            �w@        �       �                    �?0{�v��?P            @_@       �       �                   �8@,Z0R�?K             ]@        �       �                   �3@ �o_��?             9@        ������������������������       �                     @        �       �                    �?�X����?             6@        �       �                    5@      �?              @        �       �                 �{@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ���@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?؇���X�?
             ,@        ������������������������       �                     �?        �       �                    7@8�Z$���?	             *@       �       �                   �5@�C��2(�?             &@       �       �                   �4@      �?             @        ������������������������       �                      @        �       �                 ��L@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 @3�@p�C��?;            �V@        �       �                     @      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 ��@���E�?7            �U@       ������������������������       �        '             N@        �       �                    �? 7���B�?             ;@        �       �                   �<@z�G�z�?             @        ������������������������       �                      @        �       �                    ?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     6@        ������������������������       �                     "@        �       �                    @�۷E���?�            �o@        �       �                     @�q�q�?             .@       ������������������������       �                     @        �       �                    @      �?              @        ������������������������       �                     @        ������������������������       �                     @        �       �                 @3�@���KQ��?�            �m@        �       �                    �?�eP*L��?             &@       �       �                    �?�q�q�?             "@       �       �                    :@      �?              @        ������������������������       �                     �?        �       �                   �?@����X�?             @        ������������������������       �                     @        �       �                   �D@      �?             @       �       �                   �A@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       2                   �?�B�}�?�            `l@       �       �                    �?��f��?�            �j@        �       �                    �?�d�����?             3@       �       �                   �<@�r����?	             .@       �       �                     @      �?              @        �       �                 ���,@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 `v�0@r�q��?             @        ������������������������       �                     @        �       �                   �2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                     @      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �0@����H�?u            `h@        �       �                     @�q�q�?
             (@        ������������������������       �                      @        �       �                    �?���Q��?             $@        ������������������������       �                     @        �       �                 ��:@և���X�?             @       �       �                 @�%@�q�q�?             @       �       �                 pFD!@���Q��?             @       ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?               /                  �N@��GEI_�?k            �f@             ,                0��G@@`&�9�?i            �f@             	                   �?�8���?d            �e@                                @E@z�G�z�?             @                               `3@�q�q�?             @        ������������������������       �                     �?                              03�7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        
      +                   �?j���?`             e@             *                   �?BӀN��?T            �b@                                 @���g�X�?Q            `b@                              `f�)@�h����?!             L@        ������������������������       �        	             2@                                �@@�˹�m��?             C@                                 ?@؇���X�?             5@                               �*@ףp=
�?             4@                               �;@�t����?	             1@       ������������������������       �                     *@                                 =@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     1@              !                ��y @0�>���?0            �V@                                 �@@ףp=
�?             D@                             ��) @�㙢�c�?             7@                                >@P���Q�?             4@       ������������������������       �                     3@        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     1@        "      )                ���#@���J��?            �I@       #      $                  �<@ 7���B�?             ;@       ������������������������       �        	             *@        %      &                  �"@@4և���?             ,@       ������������������������       �                     &@        '      (                   ?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     8@        ������������������������       �                     @        ������������������������       �                     2@        -      .                ��?P@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        0      1                  �P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     *@        �t�bh�h*h-K ��h/��R�(KM3KK��h]�B0       �{@     �p@      L@     �f@     �F@      f@      =@      P@      @      6@      @      @              @      @                      3@      9@      E@      2@     �B@      2@      5@      &@      2@      �?      @               @      �?      @      �?                      @      $@      *@       @      *@              @       @      "@      @      @       @      @       @       @       @                       @               @      @               @      @      �?      @               @      �?      @      �?               @              @      @      @      @      @                      @      @                      0@      @      @              @      @      �?              �?      @              0@      \@      @      Q@      @      Q@             �I@      @      1@       @      *@      �?      $@              @      �?      @               @      �?      �?      �?                      �?      �?      @      �?                      @       @      @      �?              �?      @      �?       @      �?      �?      �?                      �?              �?               @       @              $@      F@      �?      1@      �?       @              @      �?      @      �?                      @              "@      "@      ;@      @      @              @      @      �?      @      �?      @                      �?       @              @      6@               @      @      ,@      �?      ,@              ,@      �?              @              &@      @               @      &@       @      &@                       @     0x@     @V@     �K@     �E@      4@      9@      (@      9@      "@       @      @       @      @      �?      @                      �?      @      �?      @                      �?       @              @      7@      @      ,@              @      @      $@      �?      $@      �?       @      �?                       @               @       @                      "@       @             �A@      2@      3@      @      @              .@      @      @      �?      �?      �?              �?      �?              @              $@      @      @              @      @      �?      @              �?      �?      @              @      �?              @              0@      *@      @      @              @      @      @               @      @      �?      �?               @      �?              �?       @              *@      @       @      @       @       @       @      �?              �?       @                      �?               @      &@      @      "@               @      @              @       @             �t@      G@      ]@      "@     �Z@      "@      2@      @      @              .@      @      @      @      �?       @      �?                       @       @      @              @       @              (@       @      �?              &@       @      $@      �?      @      �?       @              �?      �?              �?      �?              @              �?      �?              �?      �?             @V@       @      @      �?      @                      �?     �U@      �?      N@              :@      �?      @      �?       @               @      �?              �?       @              6@              "@              k@     �B@      @      $@              @      @      @              @      @             `j@      ;@      @      @      @      @      @      @      �?               @      @              @       @       @       @      �?      �?      �?      �?                      �?              �?       @             �i@      5@      h@      5@      ,@      @      *@       @      @       @      �?      �?              �?      �?              @      �?      @              �?      �?      �?                      �?      @              �?      @      �?                      @     `f@      0@       @      @       @              @      @      @              @      @       @      @       @      @      �?      @      �?                      �?      �?             `e@      (@     @e@      &@     �d@      "@      @      �?       @      �?      �?              �?      �?              �?      �?               @              d@       @     �a@       @     `a@       @     �J@      @      2@             �A@      @      2@      @      2@       @      .@       @      *@               @       @               @       @              @                      �?      1@             �U@      @      B@      @      3@      @      3@      �?      3@                      �?              @      1@              I@      �?      :@      �?      *@              *@      �?      &@               @      �?              �?       @              8@              @              2@              @       @               @      @              �?      �?              �?      �?              *@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�g?BhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMEhuh*h-K ��h/��R�(KME��h|�B@Q         p                    �?@?�p�?�           @�@               ]                   �?@�l]G���?�             p@                                   @��;�\�?q             e@                                   �?�h����?)             L@        ������������������������       �                     ;@                                   �?ܷ��?��?             =@        ������������������������       �                     @                                   �?�LQ�1	�?             7@        	       
                   �9@z�G�z�?             $@        ������������������������       �                     @                                    �?�q�q�?             @        ������������������������       �                      @                                    @      �?             @                                  <@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?                                ���`@$�q-�?	             *@       ������������������������       �                     $@                                    @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @               B                    �?h�����?H             \@              #                   �5@     ��?,             P@               "                    �?p�ݯ��?             3@                                  �?��
ц��?	             *@        ������������������������       �                     �?                                   �?�q�q�?             (@        ������������������������       �                     @                                ���@X�<ݚ�?             "@        ������������������������       �                     @                !                 @�"@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        $       =                    =@f.i��n�?            �F@       %       0                 �̌@�θ�?            �C@       &       +                   �9@���}<S�?             7@        '       (                    �?z�G�z�?             @        ������������������������       �                     �?        )       *                 pf�@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ,       /                 �Y5@�X�<ݺ?             2@       -       .                 �Y�@�8��8��?             (@        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     @        1       2                    7@     ��?             0@        ������������������������       �                     �?        3       6                    �?���Q��?             .@        4       5                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        7       <                    �?���Q��?             $@       8       ;                 @3�@z�G�z�?             @        9       :                 �?�@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        >       A                 ��y.@r�q��?             @       ?       @                 @3#%@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        C       L                    @      �?             H@        D       K                 ��T?@և���X�?	             ,@       E       J                    @���Q��?             $@       F       G                    �?z�G�z�?             @       ������������������������       �                     @        H       I                   �&@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        M       X                    �?�t����?             A@        N       S                   �;@d}h���?             ,@        O       R                   �6@�q�q�?             @       P       Q                 ��'@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        T       U                 `fv1@�C��2(�?             &@        ������������������������       �                     @        V       W                 `fV6@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        Y       \                 ��0@P���Q�?             4@        Z       [                 ��"@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             2@        ^       o                    �?�r����?8            �V@       _       h                    �?؇���X�?6             U@       `       a                    �?��2(&�?             F@        ������������������������       �                      @        b       g                 `f$@r�q��?             B@        c       d                 `fV!@؇���X�?             @        ������������������������       �                     �?        e       f                    I@r�q��?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     =@        i       j                 `f�/@R���Q�?             D@        ������������������������       �                     @        k       l                     @�X�<ݺ?             B@       ������������������������       �                     ?@        m       n                 038@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        q       �                    �?@h���?$           `|@        r       �                    �?~X�<��?3             R@       s       �                 ���<@^l��[B�?(             M@       t       �                   �=@�����H�?             B@       u       |                   @@�J�4�?             9@       v       {                   @<@@4և���?
             ,@       w       x                 ���@ףp=
�?	             $@       ������������������������       �                     @        y       z                    9@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �      �?             @        ������������������������       �                     @        }       �                    �?���!pc�?	             &@       ~                            @�q�q�?             "@        ������������������������       �                     �?        �       �                 `v�0@      �?              @       �       �                 H�Z&@z�G�z�?             @       �       �                   �<@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �2@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     &@        �       �                    @@8�A�0��?             6@       �       �                    �?�q�q�?             (@       �       �                   �8@����X�?             @        ������������������������       �                     �?        �       �                   �;@r�q��?             @        ������������������������       �                      @        �       �                    >@      �?             @       �       �                 03SA@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ��3Q@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                     �?z�G�z�?             $@       �       �                    �?      �?              @       �       �                   �I@�q�q�?             @        ������������������������       �                      @        �       �                 ��L@@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �                 Ȉ�Q@և���X�?             ,@       �       �                 =
�@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                  "&d@����X�?             @        ������������������������       �                     @        �       �                   �?@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �                       03�9@dl�"���?�            �w@       �       �                     @4?,R��?�             r@        �       �                   �M@���}<S�?)            @Q@       �       �                    �?�L#���?(            �P@       �       �                    5@Hn�.P��?$             O@        �       �                    &@؇���X�?             @        �       �                   �1@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   @A@h㱪��?             �K@       �       �                 `fF)@@-�_ .�?            �B@       ������������������������       �                     7@        �       �                   �9@؇���X�?	             ,@        ������������������������       �                      @        �       �                   �*@�q�q�?             @       �       �                    =@���Q��?             @        ������������������������       �                     �?        �       �                    @@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     2@        �       �                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �0@Ny�w��?�            `k@        �       �                     @X�<ݚ�?             "@       �       �                    �?      �?              @       �       �                 pFD!@���Q��?             @       �       �                 pf�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                 ��@�r�.kx�?�            @j@        �       �                   �;@��
ц��?             *@        �       �                 `f�@      �?              @       �       �                    6@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �                       ���#@Lvkef�?y            �h@       �       �                   �<@haLo�f�?f            �d@       �       �                    �?������?I            �^@       �       �                 �1@\#r��?H            �^@        �       �                    �?RB)��.�?            �E@       �       �                 �?$@��P���?            �D@       �       �                    �?�����H�?             B@        �       �                  s�@     ��?
             0@        ������������������������       �                     @        ������������������������       ��θ�?             *@        �       �                 ���@P���Q�?             4@        �       �                   �8@r�q��?             @        �       �                 ���@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     ,@        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?(�5�f��?.            �S@       �       �                 ��) @ �й���?+            @R@       ������������������������       �        "            �M@        �       �                 pf� @@4և���?	             ,@        ������������������������       �                     �?        ������������������������       �                     *@        �       �                    7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �                          �?      �?             F@       �       �                    �?0,Tg��?             E@        �       �                    >@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �                         �C@�d�����?             C@       �       
                  �B@��}*_��?             ;@       �       	                  @@@�q�q�?             8@       �                       ���!@b�2�tk�?
             2@       �       �                 �?�@     ��?	             0@        ������������������������       �                      @                                 �>@X�Cc�?             ,@        ������������������������       �                     @                                �?@      �?              @        ������������������������       �                     �?                              ��i @և���X�?             @                             @3�@�q�q�?             @       ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        	             &@        ������������������������       �                      @        ������������������������       �                     >@                                 @p�v>��?B            �W@                                 @z�G�z�?             @        ������������������������       �                     @                                  @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?              >                   �?@�h�|5�?>            @V@             =                   R@�4��?+            @P@             <                03�U@���h%��?*            �O@             ;                �!�N@�̚��?)            �N@             6                �TL@$��m��?$             J@             1                ��yC@���j��?             G@             0                   J@      �?             @@             #                `fF:@��
ц��?             :@              "                  �@@z�G�z�?             $@                                 �?���Q��?             @        ������������������������       �                      @               !                  �<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        $      /                  �G@      �?
             0@       %      ,                  �>@      �?	             (@       &      )                  �<@      �?              @        '      (                `fF<@      �?             @       ������������������������       �      �?              @        ������������������������       �                      @        *      +                  �B@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        -      .                �TaA@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        2      5                  �;@@4և���?	             ,@        3      4                   7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        7      8                   ;@r�q��?             @        ������������������������       �                      @        9      :                   >@      �?             @        ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                      @        ?      D                   @�8��8��?             8@       @      A                 D0T@      �?             0@       ������������������������       �                     "@        B      C                  �B@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �t�bh�h*h-K ��h/��R�(KMEKK��h]�BP       �{@     �p@     @S@     �f@     @P@     �Y@      @     �J@              ;@      @      :@              @      @      4@       @       @              @       @      @               @       @       @       @      �?       @                      �?              �?      �?      (@              $@      �?       @      �?                       @      O@      I@      :@      C@      (@      @      @      @      �?              @      @              @      @      @              @      @      �?      @                      �?      @              ,@      ?@      "@      >@       @      5@      �?      @              �?      �?      @              @      �?              �?      1@      �?      &@              @      �?      @              @      @      "@      �?              @      "@       @      @       @                      @      @      @      @      �?      �?      �?      �?                      �?      @                      @      @      �?       @      �?       @                      �?      @              B@      (@      @       @      @      @      �?      @              @      �?      �?      �?                      �?      @                      @      >@      @      &@      @      �?       @      �?      �?              �?      �?                      �?      $@      �?      @              @      �?              �?      @              3@      �?      �?      �?      �?                      �?      2@              (@     �S@      (@      R@      @      C@               @      @      >@      @      �?      �?              @      �?      @                      �?              =@      @      A@      @               @      A@              ?@       @      @              @       @                      @     �v@     �U@     �J@      3@     �F@      *@      @@      @      5@      @      *@      �?      "@      �?      @              @      �?      �?              @      �?      @               @      @      @      @              �?      @       @      @      �?      @      �?      @                      �?      �?               @      �?       @                      �?       @              &@              *@      "@      @      @       @      @      �?              �?      @               @      �?      @      �?       @               @      �?                      �?      @       @               @      @               @       @      @       @      @       @       @               @       @       @                       @       @               @               @      @      @      �?              �?      @               @      @              @       @      �?       @                      �?     �s@      Q@      o@      D@     �O@      @     �O@      @     �M@      @      @      �?       @      �?       @                      �?      @             �J@       @     �A@       @      7@              (@       @       @              @       @      @       @              �?      @      �?      �?               @      �?      �?              2@              @      �?      @                      �?               @      g@      A@      @      @      @      @      @       @      �?       @      �?                       @       @                      @      �?             �f@      =@      @      @       @      @       @      @       @                      @              @      @             �e@      7@      b@      7@     �[@      (@     �[@      (@      A@      "@      @@      "@      @@      @      *@      @      @              $@      @      3@      �?      @      �?       @      �?       @                      �?      @              ,@                      @       @              S@      @      R@      �?     �M@              *@      �?              �?      *@              @       @               @      @              �?             �@@      &@      ?@      &@      @      �?              �?      @              <@      $@      1@      $@      1@      @      &@      @      &@      @       @              "@      @      @              @      @              �?      @      @       @      @       @      �?              @      �?                       @      @                      @      &@               @              >@             �P@      <@      �?      @              @      �?      �?      �?                      �?     @P@      8@     �E@      6@     �E@      4@     �E@      2@      A@      2@     �@@      *@      4@      (@      ,@      (@       @       @      @       @       @              �?       @      �?                       @      @              @      $@      @      @      @      @      �?      @      �?      �?               @       @       @      �?              �?       @      @      �?      @                      �?              @      @              *@      �?       @      �?       @                      �?      &@              �?      @               @      �?      @      �?      �?               @      "@                       @               @      6@       @      ,@       @      "@              @       @               @      @               @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ1�.hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMEhuh*h-K ��h/��R�(KME��h|�B@Q         |                 `f�$@�6��l�?�           @�@               '                    �?�iU��2�?�            0q@               &                    �?h/��y��?0            @S@                                  �?�+e�X�?/            �R@                                   �?@�0�!��?             A@        ������������������������       �                     @                                ���@��S�ۿ?             >@        ������������������������       �                     ,@        	       
                    5@      �?
             0@        ������������������������       �                     �?                                  �<@��S�ۿ?	             .@       ������������������������       �                      @                                  �=@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @                                  �1@������?            �D@        ������������������������       �                      @               #                 `�j@��Sݭg�?            �C@              "                    �?�<ݚ�?             B@                               �Y�@4�2%ޑ�?            �A@                                   �?      �?              @                                ���@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @               !                    A@�+$�jP�?             ;@                                 �:@�q�q�?             8@        ������������������������       �                      @                                   �?�GN�z�?             6@        ������������������������       �      �?             @                                 ��(@�����H�?             2@       ������������������������       �      �?             0@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        $       %                 pF @�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        (       )                     @fhK�4�?�            �h@        ������������������������       �        
             1@        *       =                    �?Pi�b��?v            �f@        +       <                 ��i#@�P�*�?             ?@       ,       3                   �;@8�A�0��?             6@       -       2                    �?"pc�
�?             &@       .       /                 �&B@ףp=
�?             $@       ������������������������       �                     @        0       1                    4@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        4       ;                    �?���|���?             &@       5       6                 ��� @X�<ݚ�?             "@        ������������������������       �                     @        7       :                    I@z�G�z�?             @       8       9                  SE"@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@        >       C                   �0@�:pΈ��?c            �b@        ?       @                 pf�@      �?             @        ������������������������       �                     �?        A       B                 pFD!@���Q��?             @       ������������������������       �      �?             @        ������������������������       �                     �?        D       E                 @3�@      �?_             b@        ������������������������       �                      @        F       w                    �?�Z��L��?^            �a@       G       J                 ��@��IF�E�?W            �`@        H       I                 ��l@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        K       l                 @3�@�ʈD��?U             `@       L       c                 �?�@؇���X�?0            �Q@       M       \                   �;@�U�:��?'            �M@        N       [                 �1@؇���X�?             <@       O       Z                    :@�<ݚ�?             2@       P       S                 ���@      �?             0@        Q       R                 �&b@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        T       Y                   �5@$�q-�?	             *@       U       V                    4@r�q��?             @       ������������������������       �                     @        W       X                  s@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     $@        ]       b                   �@�g�y��?             ?@        ^       _                    >@�C��2(�?	             &@        ������������������������       �                     @        `       a                 �&B@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     4@        d       e                    :@�eP*L��?	             &@        ������������������������       �                     @        f       g                   �?@      �?              @        ������������������������       �                     �?        h       i                   �A@և���X�?             @        ������������������������       ��q�q�?             @        j       k                   �D@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        m       p                   �3@���#�İ?%            �M@        n       o                 ��Y @�C��2(�?             &@        ������������������������       ��q�q�?             @        ������������������������       �                      @        q       r                   �<@@��8��?             H@       ������������������������       �                     ;@        s       t                 ��)"@���N8�?             5@       ������������������������       �        
             3@        u       v                    ?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        x       {                    5@z�G�z�?             $@        y       z                    3@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        }                           @��|���?           P{@       ~       �                  x#J@
���I�?�            �s@              �                    �?������?y            `i@       �       �                    �?@��3Z��?v            �h@        �       �                     �?6uH���?&             O@        �       �                    �?�q�q�?             @       �       �                   �G@      �?             @        ������������������������       �                     �?        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�h����?!             L@       �       �                   �9@�FVQ&�?            �@@        �       �                   �7@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     9@        �       �                    6@�nkK�?             7@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     5@        �       �                    #@��5Е��?P            �`@        ������������������������       �                     $@        �       �                     �?���b��?M             _@        �       �                 `f�B@Fx$(�?              I@       �       �                 �TaA@�Q����?             D@       �       �                    �?��J�fj�?            �B@       �       �                    �?X�<ݚ�?             B@        �       �                    ?@�q�q�?             @        ������������������������       �                     �?        �       �                 ��>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �>@�eP*L��?            �@@       �       �                 ��$:@l��[B��?             =@        ������������������������       �                     @        �       �                 03k:@
j*D>�?             :@        ������������������������       �                     @        �       �                   �J@      �?             6@       �       �                   �B@�q�q�?
             .@       �       �                   @>@X�<ݚ�?             "@       �       �                 `fF<@և���X�?             @        ������������������������       �      �?             @        �       �                   �<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    H@r�q��?             @        ������������������������       �      �?             @        ������������������������       �                      @        �       �                 `fF<@؇���X�?             @        ������������������������       �                     @        �       �                   �P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        �       �                    �?������?-            �R@       �       �                    �?؇���X�?            �H@        �       �                 ���,@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?��E�B��?            �G@       �       �                   �*@�LQ�1	�?             G@       �       �                   �M@d}h���?             <@       �       �                    �?8�Z$���?             :@        ������������������������       �                      @        �       �                 `f�)@r�q��?             8@        �       �                 `f'@ףp=
�?             $@       �       �                   �5@      �?              @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                      @        �       �                   �:@d}h���?             ,@       ������������������������       �                     @        �       �                    ?@և���X�?             @        ������������������������       �                      @        �       �                   @D@z�G�z�?             @        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     2@        ������������������������       �                     �?        �       �                    :@`2U0*��?             9@        �       �                    9@ףp=
�?             $@        ������������������������       �                     @        �       �                   �E@z�G�z�?             @       �       �                   �<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     .@        ������������������������       �                     @        �       �                    �?����X�?D             \@       �       �                    �?�i�y�?(            �O@       ������������������������       �        !            �I@        �       �                     @r�q��?             (@        ������������������������       �                     �?        �       �                   �8@�C��2(�?             &@        ������������������������       �                     @        �       �                 ���`@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?`�(c�?            �H@       �       �                    �?�q�����?             9@        �       �                    �?�n_Y�K�?             *@       �       �                 @�?t@      �?              @       �       �                  �}S@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                 ��3Q@���Q��?             @        ������������������������       �                      @        �       �                 ��hU@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 `f�O@�q�q�?             (@        ������������������������       �                      @        �       �                    �?�z�G��?             $@        �       �                   �B@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �?z�G�z�?             @        ������������������������       �                     �?        �       �                 ���Y@      �?             @       ������������������������       �                     @        ������������������������       �                     �?                               03c@      �?             8@                                �?��
ц��?	             *@                                �?�<ݚ�?             "@        ������������������������       �                     @                              03�S@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     &@        	      8                   @ҐϿ<��?V            �^@       
      !                   �?X�<ݚ�?A            �V@                                 @X�Cc�?             <@        ������������������������       �                     @                                 �?�eP*L��?             6@                                �6@���!pc�?             &@        ������������������������       �                     �?                                �<@z�G�z�?             $@                                �?�<ݚ�?             "@       ������������������������       �                     @                               S�2@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?                                 �?���|���?
             &@                                 ;@      �?             @                                �2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @                                 8@և���X�?             @        ������������������������       �                      @                                �v6@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        "      #                   @f���M�?+             O@        ������������������������       �                     $@        $      %                0S�*@�θ�?&             J@        ������������������������       �                     @        &      7                �T�I@��0{9�?#            �G@       '      6                   �?�Ra����?!             F@       (      /                   �?     ��?             @@       )      .                  �8@���}<S�?             7@        *      -                   �?      �?              @        +      ,                ���0@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             .@        0      1                   )@�q�q�?             "@        ������������������������       �                     �?        2      5                   �?      �?              @        3      4                  �=@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        
             (@        ������������������������       ��q�q�?             @        9      :                   �?      �?             @@        ������������������������       �                     (@        ;      @                   �?ףp=
�?             4@        <      =                ��T?@z�G�z�?             @        ������������������������       �                     @        >      ?                   %@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        A      D                   @��S�ۿ?	             .@        B      C                   @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     (@        �t�b��>     h�h*h-K ��h/��R�(KMEKK��h]�BP       0{@     Pq@     �k@      K@     �L@      4@     �L@      2@      <@      @              @      <@       @      ,@              ,@       @              �?      ,@      �?       @              @      �?              �?      @              =@      (@               @      =@      $@      <@       @      ;@       @      @      @      �?      @      �?                      @      @              6@      @      3@      @       @              1@      @      �?      @      0@       @      ,@       @       @              @              �?              �?       @               @      �?                       @     �d@      A@      1@             `b@      A@      2@      *@      "@      *@       @      "@      �?      "@              @      �?      @      �?                      @      �?              @      @      @      @      @              �?      @      �?      �?              �?      �?                      @       @              "@              `@      5@      @      @      �?               @      @      �?      @      �?             �_@      2@               @     �_@      0@     �]@      ,@      �?       @      �?                       @     @]@      (@      N@      $@      K@      @      8@      @      ,@      @      ,@       @       @      �?       @                      �?      (@      �?      @      �?      @               @      �?       @                      �?      @                       @      $@              >@      �?      $@      �?      @              @      �?      @                      �?      4@              @      @      @              @      @              �?      @      @       @      �?      �?      @      �?       @              �?     �L@       @      $@      �?       @      �?       @             �G@      �?      ;@              4@      �?      3@              �?      �?              �?      �?               @       @      @       @      @                       @      @             �j@     �k@     �`@     �f@     �Y@     @Y@     �Y@     �W@      @     �L@       @      @       @       @              �?       @      �?       @                      �?               @      @     �J@       @      ?@       @      @              @       @                      9@      �?      6@      �?      �?              �?      �?                      5@     @X@     �B@              $@     @X@      ;@      ?@      3@      5@      3@      5@      0@      4@      0@       @      �?      �?              �?      �?      �?                      �?      2@      .@      ,@      .@      @              &@      .@              @      &@      &@      @      $@      @      @      @      @       @       @       @      �?              �?       @                       @      �?      @      �?      @               @      @      �?      @              �?      �?      �?                      �?      @              �?                      @      $@             �P@       @      E@      @      �?      �?              �?      �?             �D@      @      D@      @      6@      @      6@      @       @              4@      @      "@      �?      @      �?      �?      �?      @               @              &@      @      @              @      @               @      @      �?      @              �?      �?               @      2@              �?              8@      �?      "@      �?      @              @      �?      �?      �?      �?                      �?      @              .@                      @      @@      T@       @     �N@             �I@       @      $@      �?              �?      $@              @      �?      @              @      �?              >@      3@      (@      *@      @       @      @      @      @       @               @      @                      @       @      @               @       @      �?       @                      �?      @      @               @      @      @      @       @      @                       @      @      �?      �?              @      �?      @                      �?      2@      @      @      @      @       @      @              @       @               @      @                      @      &@              T@      E@      I@      D@      $@      2@              @      $@      (@      @       @      �?               @       @       @      @              @       @      �?       @                      �?              �?      @      @      @      �?      �?      �?      �?                      �?       @              @      @               @      @      �?      @                      �?      D@      6@              $@      D@      (@              @      D@      @     �C@      @      ;@      @      5@       @      @       @      �?       @               @      �?              @              .@              @      @              �?      @       @      �?       @      �?                       @      @              (@              �?       @      >@       @      (@              2@       @      @      �?      @              �?      �?              �?      �?              ,@      �?       @      �?              �?       @              (@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJg�)hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMGhuh*h-K ��h/��R�(KMG��h|�B�Q         |                 `f�$@<��z��?�           @�@               m                   @@@r�q��?�             p@              (                    �?����R��?�            `j@               '                    �?�\��N��?             C@                                 �9@��.k���?             A@                                  �?b�2�tk�?             2@                                 �3@j���� �?             1@                               �?@���Q��?             $@       	       
                    �?r�q��?             @        ������������������������       �                      @                                   �?      �?             @                                s�@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @                                x&�!@      �?             @       ������������������������       �                     @        ������������������������       �                     �?                                ��@؇���X�?             @                                  �5@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?               $                 �̌@     ��?             0@                                  �?�θ�?	             *@        ������������������������       �                      @                                   ;@���!pc�?             &@        ������������������������       �                      @                                ���@�q�q�?             "@        ������������������������       �                      @                !                 ���@؇���X�?             @        ������������������������       �                     @        "       #                 �&B@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        %       &                   �=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        )       ^                   �<@��D<j�?m            �e@       *       3                    �?(�����?a            `c@        +       2                   @@      �?             8@       ,       -                    5@�LQ�1	�?             7@        ������������������������       �                      @        .       1                   �7@���N8�?             5@        /       0                 ���@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     2@        ������������������������       �                     �?        4       W                    �?0�v���?R            ``@       5       6                    �?`Jj��?N             _@        ������������������������       �        
             .@        7       <                 @33@p���h�?D            @[@        8       9                     @���!pc�?             &@       ������������������������       �                     @        :       ;                    6@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        =       J                 �1@ؗp�'ʸ?=            �X@        >       ?                    7@�#-���?            �A@        ������������������������       �                     .@        @       A                   �8@R���Q�?
             4@        ������������������������       �                     �?        B       C                    :@�KM�]�?	             3@        ������������������������       �                     @        D       E                   �;@r�q��?             (@        ������������������������       �                     �?        F       G                 pf�@�C��2(�?             &@        ������������������������       �                     @        H       I                 �?$@r�q��?             @       ������������������������       �      �?             @        ������������������������       �                      @        K       L                 @3�@�i�y�?+            �O@        ������������������������       �                     4@        M       V                 ���!@ �#�Ѵ�?            �E@       N       U                   �;@`Jj��?             ?@       O       T                   �9@�t����?             1@       P       S                   �3@      �?             0@        Q       R                    2@؇���X�?             @       ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �        
             ,@        ������������������������       �                     (@        X       ]                    �?����X�?             @       Y       \                 pff@���Q��?             @       Z       [                 ���@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        _       b                    �?      �?             2@        `       a                    >@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        c       d                 �?�@և���X�?
             ,@        ������������������������       �                      @        e       h                    >@�q�q�?             (@        f       g                 ���"@      �?             @       ������������������������       �                      @        ������������������������       �                      @        i       l                 @3�@      �?              @       j       k                   �?@���Q��?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                     @        n       y                    O@=QcG��?             �G@       o       p                    �?`Ӹ����?            �F@        ������������������������       �                     @        q       r                 �?�@�7��?            �C@       ������������������������       �                     :@        s       x                    �?8�Z$���?
             *@       t       u                    �?�<ݚ�?             "@        ������������������������       �                     �?        v       w                 @3�@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        z       {                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        }       :                   @v���!��?           `|@       ~       �                     �?�!e����?�            Py@               �                   �H@����?`            @c@       �       �                  x#J@��+7��?J            �\@        �       �                   �G@D^��#��?            �D@       �       �                    �?)O���?             B@       �       �                    �?�eP*L��?            �@@        ������������������������       �                      @        �       �                    �?�P�*�?             ?@        �       �                 �ܵ<@      �?             @        ������������������������       �                      @        �       �                   �A@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    G@���Q��?             9@       �       �                   �@@\X��t�?             7@       �       �                   `@@�	j*D�?             *@        ������������������������       �                     @        ������������������������       �                     "@        �       �                    D@���Q��?             $@        ������������������������       �                     @        �       �                 `f?@�q�q�?             @       ������������������������       �      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   @C@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�x
�2�?3            �R@       ������������������������       �                     D@        �       �                    �?�!���?             A@       �       �                    �?����X�?             5@       �       �                   @D@�q�q�?             (@       �       �                    �?���!pc�?             &@        �       �                 p�w@r�q��?             @       �       �                 0c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                  "&d@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �5@�<ݚ�?             "@        ������������������������       �                     �?        �       �                 ��hU@      �?              @        �       �                 ���S@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    '@�n_Y�K�?
             *@        ������������������������       �                     @        �       �                    >@      �?             $@        ������������������������       �                     @        �       �                 03�P@����X�?             @        ������������������������       �                     @        �       �                 03�U@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                   �R@Hث3���?            �C@       �       �                    O@X�<ݚ�?             B@       �       �                    �?��S���?             >@        ������������������������       �                     &@        �       �                    �?�d�����?             3@        �       �                    �?      �?              @        ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?���|���?             &@       �       �                   �J@�z�G��?             $@        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 `f�)@�{�:��?�            `o@        �       �                   @E@��Zy�?            �C@       �       �                    �?�q�q�?            �@@       �       �                    �?� �	��?             9@       �       �                     @�8��8��?	             (@       ������������������������       �                     $@        �       �                 ��&@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�θ�?             *@        ������������������������       �                     �?        �       �                    �?r�q��?             (@       �       �                   �8@z�G�z�?             $@       �       �                    &@�q�q�?             @       �       �                   �1@���Q��?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �                          �?�ǧ\�?�            �j@        �       �                    �?`��}3��?B            �Z@       �       �                     @��C"�b�?2            �T@       �       �                    �?:ɨ��?'            �P@        �       �                    :@�t����?             1@        �       �                 ��*@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        
             *@        �       �                    �? i���t�?            �H@        �       �                 `��,@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �*@���N8�?             E@       �       �                   �;@$�q-�?             :@        ������������������������       �                     ,@        �       �                    =@r�q��?	             (@        ������������������������       �                     �?        �       �                   @D@�C��2(�?             &@        ������������������������       �                     @        �       �                   �F@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     0@        �       �                 �T)D@      �?             0@       ������������������������       �                     *@        ������������������������       ��q�q�?             @        �                          :@r�q��?             8@        �       �                     @�C��2(�?             &@        ������������������������       �                     @                                  1@      �?             @                                 @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @              
                  �B@�θ�?             *@                             `v�5@և���X�?             @        ������������������������       �                      @              	                   <@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @              '                   �?��k��?B            �Z@              $                   �?�z�G��?             I@                                �?^����?            �E@                                 �?X�Cc�?	             ,@                                P,@      �?              @        ������������������������       �                      @        ������������������������       �                     @                              03�3@      �?             @                                �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?                                  @>���Rp�?             =@                                �@@���!pc�?             &@                                �<@      �?             @                                6@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @               #                   �?�<ݚ�?             2@        !      "                ��Y.@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     (@        %      &                   �?և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        (      )                   )@>4և���?#             L@        ������������������������       �                     2@        *      3                   �?\�Uo��?             C@        +      .                0339@�E��ӭ�?
             2@        ,      -                `v�6@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        /      0                  �5@8�Z$���?             *@        ������������������������       �                     �?        1      2                   @�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        4      9                   �?ףp=
�?             4@       5      8                8#�1@؇���X�?	             ,@        6      7                   >@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     @        ;      F                   =@�q��/��?            �H@       <      =                   �?dP-���?            �G@        ������������������������       �        
             1@        >      C                ���d@�r����?             >@       ?      B                   @$�q-�?             :@        @      A                   @���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     5@        D      E                   �?      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �t�bh�h*h-K ��h/��R�(KMGKK��h]�Bp       p|@     p@     �j@     �E@     `e@      D@      4@      2@      0@      2@      &@      @      $@      @      @      @      �?      @               @      �?      @      �?      �?      �?                      �?               @      @      �?      @                      �?      @      �?      �?      �?      �?                      �?      @              �?              @      &@      @      $@               @      @       @               @      @      @       @              �?      @              @      �?      @      �?       @              �?       @      �?       @                      �?      @             �b@      6@     �a@      *@      5@      @      4@      @               @      4@      �?       @      �?              �?       @              2@              �?             @^@      $@      ]@       @      .@             @Y@       @       @      @      @              �?      @      �?                      @     @W@      @      @@      @      .@              1@      @              �?      1@       @      @              $@       @              �?      $@      �?      @              @      �?      @      �?       @             �N@       @      4@             �D@       @      =@       @      .@       @      .@      �?      @      �?      @              �?      �?      "@                      �?      ,@              (@              @       @      @       @      �?       @      �?                       @       @               @              "@      "@      @      �?              �?      @              @       @       @              @       @       @       @       @                       @       @      @       @      @               @       @      �?              @      F@      @     �E@       @      @             �B@       @      :@              &@       @      @       @      �?              @       @               @      @              @              �?      �?              �?      �?              n@     �j@     �h@      j@      I@      Z@      >@     @U@      3@      6@      3@      1@      2@      .@               @      2@      *@      @      @       @              �?      @              @      �?              .@      $@      *@      $@      "@      @              @      "@              @      @              @      @       @       @       @       @               @              �?       @               @      �?                      @      &@     �O@              D@      &@      7@      @      .@      @       @      @       @      �?      @      �?      �?              �?      �?                      @       @      @              @       @              �?               @      @      �?              �?      @      �?      @              @      �?                      @      @       @              @      @      @      @               @      @              @       @      �?       @                      �?      4@      3@      4@      0@      ,@      0@              &@      ,@      @      @      �?      @              @      �?      @                      �?      @      @      @      @      �?      @              @      �?              @                      �?      @                      @     `b@      Z@      1@      6@      &@      6@      &@      ,@      �?      &@              $@      �?      �?      �?                      �?      $@      @              �?      $@       @       @       @      @       @      @       @       @              �?       @      �?              @               @                       @      @             @`@     �T@      R@      A@     �N@      5@      G@      4@       @      .@       @       @       @                       @              *@      F@      @      @      @              @      @              D@       @      8@       @      ,@              $@       @              �?      $@      �?      @              @      �?              �?      @              0@              .@      �?      *@               @      �?      &@      *@      �?      $@              @      �?      @      �?      �?              �?      �?                       @      $@      @      @      @       @               @      @              @       @              @              M@      H@     �A@      .@      ?@      (@      "@      @      @       @               @      @              @      @       @      @              @       @              �?              6@      @       @      @      �?      @      �?      �?              �?      �?                       @      @              ,@      @       @      @       @                      @      (@              @      @              @      @              7@     �@@              2@      7@      .@      @      *@      @       @               @      @               @      &@      �?              �?      &@              &@      �?              2@       @      (@       @      �?       @               @      �?              &@              @             �E@      @     �E@      @      1@              :@      @      8@       @      @       @      @                       @      5@               @       @               @       @                       @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�]_AhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMEhuh*h-K ��h/��R�(KME��h|�B@Q                          x#J@~�Я��?�           @�@              a                    �?j;v�>��?x           ��@               Z                    @b����?t            �g@              Y                    @�q�q�?l             e@                                   @�yQ�|�?j            �d@                                   �?��.N"Ҭ?,            @Q@                                   �?�8��8��?	             (@                                    �?z�G�z�?             @        	       
                   �G@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                                  �8@0�)AU��?#            �L@                                   �?P���Q�?             4@                                 �6@�C��2(�?             &@       ������������������������       �                     @                                  �+@z�G�z�?             @       ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                    �B@               @                    �?ާb�y��?>            �W@              )                    �?�g�y��?)             O@                                03�@����X�?             <@        ������������������������       �                     @                                  �0@z�G�z�?             9@        ������������������������       �                     @               "                    �?�d�����?             3@               !                    �?      �?             @                                ��%@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        #       $                 ���@�r����?             .@        ������������������������       �                     �?        %       (                    �?@4և���?
             ,@       &       '                 pF @�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        ������������������������       �                      @        *       +                 pf�@ҳ�wY;�?             A@        ������������������������       �                     @        ,       -                    7@>���Rp�?             =@        ������������������������       �                     @        .       7                    �?8����?             7@       /       2                   �;@�θ�?	             *@        0       1                   �9@      �?             @        ������������������������       �                      @        ������������������������       �                      @        3       4                 `�X!@�����H�?             "@       ������������������������       �                     @        5       6                  SE"@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        8       ?                   �=@���Q��?             $@       9       :                 pf�'@և���X�?             @        ������������������������       �                     �?        ;       >                    ;@�q�q�?             @       <       =                 @3�/@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        A       N                    �?����e��?            �@@       B       M                 �A7@      �?             0@       C       H                 P��%@z�G�z�?
             .@        D       E                    $@      �?             @        ������������������������       �                     �?        F       G                   �7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        I       J                    0@�C��2(�?             &@       ������������������������       �                     @        K       L                 03S1@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        O       X                 `v�6@��.k���?
             1@       P       Q                 ��"@���!pc�?             &@        ������������������������       �                     �?        R       W                    �?z�G�z�?             $@       S       V                 ���.@����X�?             @        T       U                   �<@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        [       `                   �>@��s����?             5@       \       ]                    @�X�<ݺ?             2@       ������������������������       �                     *@        ^       _                 ���3@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        b       �                     �?�#߆;s�?            z@        c       d                   �;@������?%             Q@        ������������������������       �                     @        e       l                    �?     ��?$             P@        f       k                    �?�8��8��?             (@       g       h                 ��L@@؇���X�?             @       ������������������������       �                     @        i       j                   �B@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        m       �                    �? s�n_Y�?             J@       n                           R@�q�q��?             H@       o       ~                    K@�3Ea�$�?             G@       p       }                   �H@�������?             A@       q       x                 `f�;@     ��?             @@       r       s                   �9@և���X�?             ,@        ������������������������       �                     @        t       w                   �E@      �?              @       u       v                   �?@r�q��?             @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �      �?              @        y       |                   �<@�X�<ݺ?	             2@       z       {                   �>@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     (@        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?��Mjs�?�            �u@       �       �                    �?�r����?�            �q@       �       �                     @h�Q�j��?�            �q@        �       �                    @@�����?,            �R@       �       �                    �?8�Z$���?            �C@        �       �                   �9@      �?             @        ������������������������       �                     �?        �       �                    =@���Q��?             @       �       �                 ���,@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�C��2(�?            �@@       �       �                    5@HP�s��?             9@        �       �                   �1@      �?             @        ������������������������       �                      @        �       �                   �'@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �;@���N8�?             5@       ������������������������       �                     &@        �       �                    =@ףp=
�?             $@       �       �                    @�����H�?             "@       ������������������������       �                     @        �       �                   �*@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �7@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?��?^�k�?            �A@        ������������������������       �                      @        �       �                 `f'@Pa�	�?            �@@        �       �                   �P@z�G�z�?             @       �       �                   @H@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     <@        �       �                 ��@�����?�            �i@        �       �                    �?     ��?             0@       �       �                    �?�q�q�?
             .@        ������������������������       �                     @        �       �                 ���@�eP*L��?             &@       �       �                 ���	@؇���X�?             @        �       �                    6@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?��K�# �?{            �g@        �       �                  ��@�iʫ{�?"            �J@        �       �                   �6@ �q�q�?             8@        ������������������������       �                     �?        ������������������������       �                     7@        �       �                    �?�c�Α�?             =@       �       �                    �?R�}e�.�?             :@        �       �                 @3s+@�q�q�?             "@       �       �                 �� @؇���X�?             @       �       �                    ?@z�G�z�?             @        �       �                   �<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                 ��(@������?
             1@       �       �                   �<@����X�?             ,@       ������������������������       �                      @        �       �                   �>@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                 �*@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ��@�q��/��?Y            @a@        ������������������������       �                     3@        �       �                    �?��5Վ3�?L            �]@       �       �                   �<@���AS��?F            @[@       �       �                 �1@ףp=
�?/            �Q@        �       �                 �?$@�q�q�?             @        ������������������������       �                      @        �       �                   �6@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                 �?�@     p�?+             P@        ������������������������       �                     4@        �       �                 @�!@�Ra����?             F@       �       �                 ��) @д>��C�?             =@       �       �                   �3@��2(&�?             6@        ������������������������       �                     @        ������������������������       �                     3@        �       �                 ��i @����X�?             @        ������������������������       �                     �?        �       �                 pf� @r�q��?             @        ������������������������       �                      @        �       �                    8@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             .@        �       �                   �=@:�&���?            �C@        ������������������������       �                     @        �       �                   �F@�����H�?             B@       �       �                   �@؇���X�?             <@        ������������������������       �                     �?        �       �                   �E@�����H�?             ;@       �       �                 @3�@ �q�q�?             8@        �       �                 �?�@�����H�?             "@        ������������������������       �                     @        �       �                   �A@r�q��?             @       ������������������������       �      �?             @        ������������������������       �                      @        ������������������������       �        	             .@        �       �                 @3�@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 �&B@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        �       �                 ���/@      �?             @       ������������������������       �                      @        ������������������������       �                      @                                  @R=6�z�?*            @P@                                '@^n����?)             N@                                 @4���C�?            �@@        ������������������������       �                     @                                  @|��?���?             ;@        ������������������������       �                     $@                                 @@�0�!��?
             1@                                 �?�q�q�?             "@       ������������������������       �                     @        	      
                pf�C@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     ;@        ������������������������       �                     @              >                   �?lwY���?B            @Z@             1                 "�`@r�q��?6             U@             ,                    @�����H�?)            �O@             '                ���X@x�}b~|�?&            �L@             &                    �?���.�6�?             G@                               �5@t��ճC�?             F@                              ��gS@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?              %                   �?���N8�?             E@                             @3�L@�FVQ&�?            �@@                                 �?r�q��?             @        ������������������������       �                     �?                                @K@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?                                  �? 7���B�?             ;@       ������������������������       �                     6@        !      "                  @B@z�G�z�?             @        ������������������������       �                      @        #      $                  �G@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                      @        (      +                pf�Z@"pc�
�?             &@        )      *                   D@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        -      .                   ;@�q�q�?             @        ������������������������       �                     @        /      0                   >@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        2      7                  �<@�q�q�?             5@        3      6                   4@      �?              @        4      5                   $@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        8      =                ���f@$�q-�?             *@        9      :                   �?      �?             @        ������������������������       �                      @        ;      <                   H@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        ?      D                   �?؇���X�?             5@        @      A                   �?�q�q�?             "@        ������������������������       �                     �?        B      C                   :@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     (@        �t�bh�h*h-K ��h/��R�(KMEKK��h]�BP       �{@     �p@     �y@     �h@     �P@     �^@     �H@     �]@     �F@     �]@       @     �P@      �?      &@      �?      @      �?      �?              �?      �?                      @              @      �?      L@      �?      3@      �?      $@              @      �?      @      �?       @               @              "@             �B@     �E@      J@      >@      @@       @      4@      @              @      4@              @      @      ,@      @      �?      �?      �?              �?      �?               @               @      *@      �?              �?      *@      �?      &@              &@      �?                       @      6@      (@              @      6@      @      @              0@      @      $@      @       @       @       @                       @       @      �?      @              �?      �?              �?      �?              @      @      @      @      �?               @      @       @      �?              �?       @                      @      @              *@      4@      @      (@      @      (@       @       @      �?              �?       @               @      �?              �?      $@              @      �?      @      �?                      @      �?              "@       @      @       @      �?               @       @       @      @       @       @       @                       @              @              @      @              @              1@      @      1@      �?      *@              @      �?              �?      @                      @     �u@     @R@      J@      0@              @      J@      (@      &@      �?      @      �?      @               @      �?              �?       @              @             �D@      &@     �B@      &@     �B@      "@      9@      "@      9@      @       @      @      @               @      @      �?      @      �?       @              @      �?      �?      1@      �?      "@      �?              �?      "@               @                       @      (@                       @      @             Pr@     �L@     �n@      C@     �n@      B@     �P@      @     �@@      @      @      @      �?               @      @      �?      @              @      �?              �?              >@      @      7@       @      @      �?       @              �?      �?              �?      �?              4@      �?      &@              "@      �?       @      �?      @              �?      �?              �?      �?              �?              @      �?      @                      �?      A@      �?       @              @@      �?      @      �?      �?      �?      �?                      �?      @              <@             @f@      =@      &@      @      $@      @      @              @      @      @      �?      �?      �?      �?                      �?      @                      @      �?             �d@      8@      F@      "@      7@      �?              �?      7@              5@       @      3@      @      @      @      @      �?      @      �?      �?      �?      �?                      �?      @               @                       @      *@      @      $@      @       @               @      @              @       @              @               @      �?              �?       @             �^@      .@      3@              Z@      .@     �W@      ,@     �O@      @      @       @       @               @       @               @       @             �M@      @      4@             �C@      @      8@      @      3@      @              @      3@              @       @              �?      @      �?       @              @      �?      @                      �?      .@              @@      @              @      @@      @      8@      @              �?      8@      @      7@      �?       @      �?      @              @      �?      @      �?       @              .@              �?       @               @      �?               @              "@      �?              �?      "@               @       @       @                       @      G@      3@     �D@      3@      ,@      3@              @      ,@      *@              $@      ,@      @      @      @      @               @      @              @       @               @              ;@              @              @@     @R@      ,@     �Q@      @      L@      @      J@      @     �E@      @     �D@      �?      �?      �?                      �?       @      D@       @      ?@      �?      @              �?      �?      @              @      �?              �?      :@              6@      �?      @               @      �?       @      �?                       @              "@               @       @      "@       @      �?              �?       @                       @       @      @              @       @      �?       @                      �?      @      ,@      @       @      �?       @      �?                       @      @              �?      (@      �?      @               @      �?      �?      �?                      �?              "@      2@      @      @      @              �?      @       @               @      @              (@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJL�OhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMmhuh*h-K ��h/��R�(KMm��h|�B@[         �                     @������?�           @�@               [                    �?����e��?�            �s@                                  �?䖪@���?�            �g@                                  �H@��ɉ�?/            @P@                                   �? �Jj�G�?'            �K@        ������������������������       �                     :@                                   �?XB���?             =@              	                 `f�)@�}�+r��?             3@        ������������������������       �                     @        
                        ��*@�8��8��?
             (@                                  :@      �?              @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@                                  @J@ףp=
�?             $@                                   �?�q�q�?             @                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @               :                 ��=@� ��1�?V            �^@                                  �?�Zl�i��?4            @T@        ������������������������       �                     @               /                 ��$:@�KM�]�?1             S@              .                   �*@85�}C�?(            �N@                                  @X�EQ]N�?            �E@        ������������������������       �                     @               %                   �C@4?,R��?             B@                                `fF)@h�����?             <@        ������������������������       �                     .@        !       "                   �:@$�q-�?	             *@       ������������������������       �                     &@        #       $                    =@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        &       )                 `f'@      �?              @        '       (                   �P@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        *       +                 `f�)@���Q��?             @        ������������������������       �                     �?        ,       -                    G@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     2@        0       1                 03k:@z�G�z�?	             .@        ������������������������       �                     �?        2       9                 `f�;@؇���X�?             ,@       3       8                   @L@r�q��?             (@       4       7                    H@����X�?             @       5       6                   @B@r�q��?             @        ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ;       P                 0�&C@�ՙ/�?"             E@        <       O                   �A@r�q��?             8@       =       F                   @A@D�n�3�?             3@       >       ?                   �;@���Q��?             $@        ������������������������       �                     �?        @       A                    �?X�<ݚ�?             "@        ������������������������       �                      @        B       E                   �>@և���X�?             @       C       D                   �<@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        G       H                 ���=@�<ݚ�?             "@        ������������������������       �                      @        I       N                   �P@����X�?             @       J       M                   �J@r�q��?             @       K       L                   �H@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        Q       Z                 p�w@r�q��?             2@       R       S                    *@�t����?             1@        ������������������������       �                     �?        T       Y                   �;@      �?             0@        U       X                    �?�q�q�?             @       V       W                 ���Z@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     *@        ������������������������       �                     �?        \       �                    �?������?N             `@       ]       p                     �?���>4��?1             U@       ^       o                   @I@�\�u��?            �I@       _       n                    �?���|���?             F@       `       m                   �H@8�$�>�?            �E@       a       l                   �G@�d�����?             C@       b       k                    D@�4�����?             ?@       c       d                    �?      �?             <@        ������������������������       �                     .@        e       j                   �B@��
ц��?	             *@       f       i                 `f�N@�q�q�?             (@        g       h                 `fFJ@      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        q       �                    @@:ɨ��?            �@@       r       y                    9@�G�z��?             4@        s       x                     @�<ݚ�?             "@       t       w                    �?      �?              @        u       v                 ��m1@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        z                           �?���|���?             &@       {       ~                    ;@�<ݚ�?             "@        |       }                    6@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                   �7@$�q-�?             *@        ������������������������       �                     @        �       �                    �?ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        �       �                    :@f.i��n�?            �F@        ������������������������       �                     $@        �       �                    H@���Q��?            �A@       �       �                   �8@8^s]e�?             =@        �       �                    �?8�Z$���?	             *@       �       �                    @����X�?             @        ������������������������       �                     �?        �       �                   pI@r�q��?             @       �       �                    �?�q�q�?             @        ������������������������       �                     �?        �       �                    +@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?     ��?             0@       �       �                    <@      �?              @        �       �                    �?      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                 Ј2T@      �?              @       �       �                    �?r�q��?             @        ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                 03�S@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?>b3C[
�?�            �x@        �       �                 `v�6@�7i���?A            �Y@       �       �                   �:@gO�~k�?4            @T@       �       �                  s�@v ��?            �E@        ������������������������       �                     @        �       �                 @33"@X�<ݚ�?             B@        �       �                 @� @�z�G��?             4@       �       �                    @���Q��?	             .@       �       �                    �?X�Cc�?             ,@       �       �                 ���@�n_Y�K�?             *@       �       �                    �?�q�q�?             (@        ������������������������       �                     �?        �       �                 pff@���|���?             &@       �       �                    4@�q�q�?             "@        ������������������������       �                     @        �       �                   �7@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                   �8@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?      �?             0@        �       �                    9@����X�?             @       �       �                    �?���Q��?             @        ������������������������       �                     �?        �       �                    �?      �?             @        �       �                    4@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    6@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�����H�?             "@       �       �                    �?؇���X�?             @        ������������������������       �                     �?        �       �                 pf�0@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 �̌@�I�w�"�?             C@        �       �                  s�@��S�ۿ?             .@        ������������������������       �                      @        �       �                    �?$�q-�?             *@       ������������������������       �                     (@        ������������������������       �                     �?        �       �                   @B@�LQ�1	�?             7@       �       �                    @�X����?             6@       �       �                    @@����X�?             5@       �       �                 �?�@�q�q�?             2@        ������������������������       �                     �?        �       �                    �?�t����?
             1@        �       �                    �?؇���X�?             @       �       �                   �<@z�G�z�?             @       �       �                  S�2@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �;@���Q��?             $@        ������������������������       �                      @        �       �                    �?      �?              @       �       �                    �?և���X�?             @        �       �                 ��� @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ��1@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    @؇���X�?             5@        ������������������������       �                     @        ������������������������       �                     2@        �       �                   �	@��S�U�?�            Pr@        �       �                   �>@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       R                   �?,&1��?�            r@       �       �                    !@�K��E/�?�            �k@        ������������������������       �                     @        �       /                  �<@������?�            @k@       �       
                   �?@݈g>h�?_             c@        �                       ��*@H%u��?             9@       �                        ���@���}<S�?             7@        ������������������������       �                     @                                @@      �?             0@                                9@"pc�
�?             &@        ������������������������       �                     �?                                @<@z�G�z�?             $@       ������������������������       ��<ݚ�?             "@        ������������������������       �                     �?        ������������������������       �                     @              	                  �2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                              ��@4Jı@�?R            �_@                                 7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                �0@Ȓ�g;�?P             _@                              pFD!@z�G�z�?             $@                             pf�@����X�?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     @              ,                �!&B@Xl���?L            �\@                             ��@ ��WV�?H             Z@        ������������������������       �                     6@                                 �?������?8            �T@        ������������������������       �                     �?              !                �1@H�!b	�?7            @T@                              �?$@"pc�
�?             &@                                 ;@z�G�z�?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @                                 �6@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        "      '                  �3@��?^�k�?1            �Q@        #      &                ��Y @�C��2(�?             &@        $      %                �?�@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        (      )                  �:@P����?)            �M@        ������������������������       �                     ?@        *      +                  �;@h�����?             <@        ������������������������       �                     �?        ������������������������       �                     ;@        -      .                   ;@�z�G��?             $@        ������������������������       �                     �?        ������������������������       ��<ݚ�?             "@        0      9                �&B@"pc�
�?*            �P@        1      2                ��}@�nkK�?             7@       ������������������������       �        	             *@        3      8                ��@ףp=
�?             $@       4      7                   �?؇���X�?             @       5      6                   >@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        :      M                ��i @�%^�?            �E@       ;      B                �?�@�4�����?             ?@        <      A                  @@@������?             1@        =      >                  �=@�q�q�?             @        ������������������������       �                      @        ?      @                   ?@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     &@        C      J                  @B@և���X�?	             ,@       D      I                  �@@�z�G��?             $@       E      F                   ?@      �?             @        ������������������������       �                     �?        G      H                @3�@���Q��?             @       ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        K      L                  �D@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        N      O                ���"@�8��8��?	             (@       ������������������������       �                     $@        P      Q                   (@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        S      f                  �9@�����?,             Q@       T      _                   3@V������?            �B@       U      Z                   @�������?             >@        V      W                ��|2@      �?             @        ������������������������       �                     �?        X      Y                   �?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        [      ^                   @r�q��?             8@       \      ]                   +@���|���?             &@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     *@        `      a                   6@և���X�?             @        ������������������������       �                      @        b      c                  �8@���Q��?             @        ������������������������       �                      @        d      e                (3�)@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        g      h                   �?`Jj��?             ?@       ������������������������       �                     1@        i      j                 �v6@؇���X�?             ,@        ������������������������       �                     "@        k      l                   �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �t�b�      h�h*h-K ��h/��R�(KMmKK��h]�B�        |@     `p@     @c@     `d@     @Y@     �U@       @     �O@      �?      K@              :@      �?      <@      �?      2@              @      �?      &@      �?      @      �?       @              @              @              $@      �?      "@      �?       @      �?      �?      �?                      �?              �?              @     �X@      8@     @R@       @      @              Q@       @      L@      @      C@      @      @              ?@      @      ;@      �?      .@              (@      �?      &@              �?      �?              �?      �?              @      @      �?       @               @      �?              @       @      �?               @       @               @       @              2@              (@      @              �?      (@       @      $@       @      @       @      @      �?      @               @      �?              �?      @               @              :@      0@      &@      *@      &@       @      @      @              �?      @      @               @      @      @      �?      @              @      �?              @              @       @       @              @       @      @      �?       @      �?       @                      �?      @                      �?              @      .@      @      .@       @              �?      .@      �?       @      �?      �?      �?              �?      �?              �?              *@                      �?     �J@      S@     �C@     �F@      0@     �A@      0@      <@      .@      <@      $@      <@      $@      5@      @      5@              .@      @      @      @      @      @      @      @                      @      @                      �?      @                      @      @              �?                      @      7@      $@      &@      "@      @       @      @      �?       @      �?              �?       @              @                      �?      @      @       @      @       @       @               @       @                      @       @              (@      �?      @              "@      �?              �?      "@              ,@      ?@              $@      ,@      5@      "@      4@       @      &@       @      @      �?              �?      @      �?       @              �?      �?      �?              �?      �?                      @              @      @      "@       @      @       @       @               @       @                      @      @      @      @      �?      @               @      �?              �?       @                       @      @      �?              �?      @             �r@     �X@     �G@     �K@      =@      J@      4@      7@              @      4@      0@      ,@      @      "@      @      "@      @       @      @       @      @      �?              @      @      @      @      @               @      @              @       @              �?      �?      �?                      �?              �?      �?                      �?      @              @      $@      @       @      @       @      �?               @       @      �?      �?              �?      �?              �?      �?      �?                      �?       @              �?       @      �?      @              �?      �?      @              @      �?                       @      "@      =@      �?      ,@               @      �?      (@              (@      �?               @      .@      @      .@      @      .@      @      (@      �?              @      (@      �?      @      �?      @      �?       @      �?                       @               @               @      @      @               @      @      @      @      @      �?      �?      �?                      �?       @      @              @       @              �?                      @      �?              �?              2@      @              @      2@              o@      F@       @       @               @       @             �n@      E@      h@      =@              @      h@      :@     @a@      ,@      6@      @      5@       @      @              ,@       @      "@       @      �?               @       @      @       @      �?              @              �?      �?      �?                      �?      ]@      &@      �?       @      �?                       @     �\@      "@       @       @      @       @      �?              @       @      @             �Z@      @      Y@      @      6@             �S@      @      �?             @S@      @      "@       @      @      �?       @               @      �?      @      �?              �?      @              Q@       @      $@      �?      @      �?      @                      �?      @              M@      �?      ?@              ;@      �?              �?      ;@              @      @              �?      @       @      K@      (@      6@      �?      *@              "@      �?      @      �?      @      �?              �?      @              @              @              @@      &@      5@      $@      *@      @       @      @               @       @       @       @                       @      &@               @      @      @      @      @      @      �?               @      @       @      �?               @      @              �?      @      �?       @              �?      &@      �?      $@              �?      �?              �?      �?             �K@      *@      :@      &@      7@      @      @      @              �?      @       @      @                       @      4@      @      @      @              @      @              *@              @      @               @      @       @       @              �?       @               @      �?              =@       @      1@              (@       @      "@              @       @               @      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ��lhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM#huh*h-K ��h/��R�(KM#��h|�B�H         l                     @4�<����?�           @�@                                   �?x����?�            �r@                                    �?���f�?Y             `@               	                    �?�X�<ݺ?'             K@                                  �H@ ��WV�?             :@       ������������������������       �                     4@                                  �J@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        
                        ���a@@4և���?             <@       ������������������������       �                     7@                                   ;@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @                                   �?��
���?2            �R@                                 �;@�nkK�?             G@                                  �6@�r����?             .@        ������������������������       �                     @                                ��m1@�<ݚ�?             "@                               ���*@؇���X�?             @                                 �'@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �      �?             @        ������������������������       �                      @                                  �9@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ?@        ������������������������       �                     =@                                   (@x���@O�?o             e@        ������������������������       �                     "@                U                     �?��Q���?h             d@       !       0                 ��=@��+7��?:             W@        "       #                    �?$�q-�?             :@        ������������������������       �                     @        $       )                 03k:@ףp=
�?             4@        %       &                   �D@z�G�z�?             @        ������������������������       �                     @        '       (                   �9@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        *       /                    J@��S�ۿ?             .@        +       .                 `f�;@r�q��?             @       ,       -                   @G@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        1       H                   �B@�q�q�?,            �P@       2       G                    �?�s��:��?             C@       3       4                   �8@�q�q�?             B@        ������������������������       �                     @        5       :                    �?�g�y��?             ?@        6       9                 �D�G@�q�q�?             (@        7       8                 `f�A@      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ;       @                    �?D�n�3�?             3@       <       ?                 ��yC@      �?             $@       =       >                   @>@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        A       F                   @B@�q�q�?             "@       B       C                   @K@؇���X�?             @        ������������������������       �                     @        D       E                 `f�N@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        I       T                    �?�>4և��?             <@       J       O                    �?ȵHPS!�?             :@       K       N                    @@8�Z$���?	             *@        L       M                   �J@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        P       S                 p"�S@$�q-�?             *@        Q       R                 �UwR@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        V       c                   �<@����p�?.             Q@        W       ^                 ��\+@؇���X�?             <@       X       ]                    5@�����?             5@        Y       Z                   �2@�<ݚ�?             "@        ������������������������       �                     @        [       \                   �'@�q�q�?             @       ������������������������       �      �?             @        ������������������������       �                      @        ������������������������       �        
             (@        _       b                    �?����X�?             @       `       a                 `��,@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        d       k                   @A@�(\����?             D@        e       f                    �?P���Q�?             4@        ������������������������       �                     @        g       j                    �?@4և���?             ,@       h       i                   �@@      �?              @        ������������������������       �                     �?        ������������������������       �؇���X�?             @        ������������������������       �                     @        ������������������������       �                     4@        m       n                    �?�G�5��?�            �y@        ������������������������       �                     @        o                       @3�4@������?�            �y@       p       �                    �?�y�o%[�?�            pt@       q       ~                   �0@^�g��?�            pp@        r       w                    �?r�q��?             8@        s       v                    �?ףp=
�?             $@        t       u                    @      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        x       y                    .@����X�?             ,@        ������������������������       �                     @        z       {                 pf�@X�<ݚ�?             "@        ������������������������       �                      @        |       }                 pFD!@և���X�?             @        ������������������������       �z�G�z�?             @        ������������������������       �                      @               �                    �?^wUBO��?�            �m@        �       �                 `f�%@l��[B��?%             M@       �       �                    �?� �	��?             I@       �       �                    �?Tt�ó��?            �H@        �       �                    4@�ՙ/�?             5@        ������������������������       �                      @        �       �                 pF @�����?             3@       �       �                    �?������?             1@        ������������������������       �                     �?        �       �                 ���@      �?
             0@        ������������������������       �                     @        �       �                 ���@$�q-�?	             *@        ������������������������       �                     @        �       �                    9@ףp=
�?             $@        ������������������������       �                      @        �       �                 �&B@      �?              @       ������������������������       �؇���X�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ��}@��X��?             <@        ������������������������       �                      @        �       �                   �;@R�}e�.�?             :@       �       �                    �?p�ݯ��?             3@       �       �                   �9@�q�q�?             2@       �       �                  �#@؇���X�?             ,@       �       �                   �6@�C��2(�?             &@       �       �                  p @r�q��?             @        �       �                    4@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 �[$@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?      �?              @        ������������������������       �                     @        �       �                    �?���Q��?             @        ������������������������       �                     �?        �       �                 �a*@      �?             @        ������������������������       �                     �?        �       �                    @�q�q�?             @       �       �                   �<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?��CC`)�?u            �f@        �       �                 @3s+@�8��8��?             8@       �       �                 ���@�nkK�?             7@        ������������������������       �                     "@        �       �                   @@@4և���?             ,@       �       �                    9@�����H�?             "@        ������������������������       �                     �?        �       �                    =@      �?              @       ������������������������       �؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �:@�Z��=��?b            �c@        �       �                 �?$@�nkK�?             G@        ������������������������       �                     2@        �       �                 ��L@@4և���?             <@        �       �                   �6@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 �?�@`2U0*��?             9@        ������������������������       �                     *@        �       �                   �3@�8��8��?	             (@       �       �                 ��Y @؇���X�?             @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�ȼB���?E            �[@        �       �                    >@z�G�z�?             4@       �       �                   �<@������?             1@       �       �                 ��(@     ��?
             0@       �       �                  s�@      �?             (@        ������������������������       �                     @        ������������������������       ��q�q�?             "@        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?H�g�}N�?7            �V@       �       �                   �;@��2(&�?4             V@        ������������������������       �                     @        �       �                   �<@�����?1             U@        �       �                 ��) @ qP��B�?            �E@       ������������������������       �                    �A@        �       �                 pf� @      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ���"@��r._�?            �D@       �       �                 �&B@������?            �B@        ������������������������       �                     0@        �       �                   �@��s����?             5@        ������������������������       �                      @        �       �                 �?�@�KM�]�?             3@        ������������������������       �                     @        �       �                 @3�@r�q��?             (@        ������������������������       �                     �?        �       �                 ��!@�C��2(�?             &@       �       �                   �@@      �?              @       �       �                    ?@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    ?@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �                          @     ��?*             P@       �       �                    .@���Q��?(             N@        �       �                    �?��2(&�?             6@       �       �                 P�@r�q��?             2@        ������������������������       �                     @        �       �                   �*@      �?
             (@        ������������������������       �                      @        �       �                 pff!@ףp=
�?             $@        �       �                   �6@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �                       03;4@�s��:��?             C@                                 +@�'�=z��?            �@@        ������������������������       �                     @                                 �?*;L]n�?             >@                                �?      �?             :@                                �?������?	             1@        ������������������������       �                     @              	                   ;@�q�q�?             (@                                 9@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        
                      03�1@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @                                 @ wVX(6�?,            @T@                                 @�+$�jP�?
             ;@       ������������������������       �                     2@                                 @X�<ݚ�?             "@        ������������������������       �                     @                                 @z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?              "                   �? 7���B�?"             K@              !                    @8�Z$���?             *@                                ;@"pc�
�?             &@        ������������������������       �                     �?                              �T)D@ףp=
�?             $@        ������������������������       �                     @                                  >@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                    �D@        �t�bh�h*h-K ��h/��R�(KM#KK��h]�B0        |@     �p@      a@     @d@      @      _@      @     �I@      �?      9@              4@      �?      @      �?                      @       @      :@              7@       @      @       @                      @       @     @R@       @      F@       @      *@              @       @      @      �?      @      �?      @              �?      �?      @               @      �?      �?              �?      �?                      ?@              =@     ``@      C@              "@     ``@      =@      Q@      8@      8@       @      @              2@       @      @      �?      @              �?      �?      �?                      �?      ,@      �?      @      �?       @      �?       @                      �?      @              "@              F@      6@      5@      1@      5@      .@      @              0@      .@      @      @      @      @              @      @                      @      &@       @      @      @       @      @       @                      @      @              @      @      @      �?      @               @      �?              �?       @                       @               @      7@      @      7@      @      &@       @      �?       @               @      �?              $@              (@      �?      @      �?      @                      �?       @                       @     �O@      @      8@      @      3@       @      @       @      @              @       @       @       @       @              (@              @       @      @       @               @      @               @             �C@      �?      3@      �?      @              *@      �?      @      �?      �?              @      �?      @              4@             �s@     �Y@              @     �s@      X@     �m@     @V@     @i@     �N@      &@      *@      �?      "@      �?      @              @      �?                      @      $@      @      @              @      @       @              @      @      �?      @       @             �g@      H@      >@      <@      <@      6@      ;@      6@       @      *@       @              @      *@      @      *@              �?      @      (@      @              �?      (@              @      �?      "@               @      �?      @      �?      @              �?       @              3@      "@               @      3@      @      (@      @      (@      @      (@       @      $@      �?      @      �?       @      �?       @                      �?      @              @               @      �?              �?       @                      @              �?      @              �?               @      @              @       @      @      �?              �?      @              �?      �?       @      �?      �?      �?                      �?              �?      d@      4@      6@       @      6@      �?      "@              *@      �?       @      �?      �?              @      �?      @      �?      �?              @                      �?     `a@      2@      F@       @      2@              :@       @       @      �?              �?       @              8@      �?      *@              &@      �?      @      �?      �?      �?      @              @             �W@      0@      0@      @      *@      @      *@      @      "@      @      @              @      @      @                      �?      @             �S@      (@      S@      (@              @      S@       @      E@      �?     �A@              @      �?              �?      @              A@      @     �@@      @      0@              1@      @               @      1@       @      @              $@       @              �?      $@      �?      @      �?      @      �?      @                      �?      @              @              �?      @              @      �?              @              B@      <@      B@      8@      3@      @      .@      @      @              "@      @               @      "@      �?      �?      �?              �?      �?               @              @              1@      5@      1@      0@              @      1@      *@      *@      *@      @      *@              @      @       @       @      �?              �?       @               @      @              @       @              "@              @                      @              @     �R@      @      6@      @      2@              @      @              @      @      �?      @                      �?      J@       @      &@       @      "@       @              �?      "@      �?      @              @      �?      @                      �?       @             �D@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�-#hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM5huh*h-K ��h/��R�(KM5��h|�B@M         �                     @4�<����?�           @�@                                  �'@�!�����?�            pt@                                   @д>��C�?             =@        ������������������������       �        	             &@                                  �E@�E��ӭ�?             2@                                  &@d}h���?	             ,@                                 �;@�θ�?             *@               	                    �?և���X�?             @        ������������������������       �                      @        
                          �5@z�G�z�?             @                                 �1@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?                                   N@      �?             @        ������������������������       �                      @        ������������������������       �                      @               }                 �D�O@ўKr��?�            �r@              p                    �?<�����?x            �i@              '                    �?���t���?l            �g@               &                    �?x�}b~|�?"            �L@                                   �?�*/�8V�?            �G@                                   �?�z�G��?             $@                                   �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @               %                   �;@@-�_ .�?            �B@                                    �?"pc�
�?             &@        ������������������������       �                     @        !       $                   �9@�q�q�?             @       "       #                   �3@z�G�z�?             @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     :@        ������������������������       �                     $@        (       )                    +@ތux��?J            ``@        ������������������������       �                     @        *       O                     �?�w��@�?F            �_@        +       L                    �?�T��5m�?"            �P@       ,       I                    �?Z��Yo��?             O@       -       4                    �?l`N���?            �J@        .       3                   �L@X�<ݚ�?             "@       /       0                 �ܵ<@�q�q�?             @        ������������������������       �                     �?        1       2                 `f�B@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        5       H                   �>@8�A�0��?             F@       6       7                   �;@��.k���?             A@        ������������������������       �                     @        8       A                   @=@և���X�?             <@       9       :                   �9@      �?	             0@        ������������������������       �                      @        ;       <                 03k:@����X�?             ,@        ������������������������       �                     �?        =       >                   `G@�θ�?             *@        ������������������������       �                      @        ?       @                   �K@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        B       C                   �<@�q�q�?             (@        ������������������������       �                     @        D       G                   @>@      �?              @       E       F                   @K@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     $@        J       K                    �?�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        M       N                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        P       g                    �?(2��R�?$            �M@       Q       X                    �?     ��?             @@        R       W                    �?r�q��?             @       S       T                   �9@z�G�z�?             @        ������������������������       �                      @        U       V                 ���,@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        Y       f                   �*@���B���?             :@       Z       [                 `f�)@      �?             4@        ������������������������       �                     �?        \       ]                   �;@�d�����?             3@        ������������������������       �                     $@        ^       _                    =@X�<ݚ�?             "@        ������������������������       �                      @        `       e                   @D@և���X�?             @       a       b                    @@z�G�z�?             @        ������������������������       �                     �?        c       d                   @B@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        h       i                    �?�>����?             ;@        ������������������������       �                     @        j       o                    �?ףp=
�?             4@       k       n                   �@@r�q��?             (@        l       m                   �<@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        q       r                   �7@�d�����?             3@        ������������������������       �                      @        s       v                    �?�eP*L��?             &@        t       u                   `A@      �?             @        ������������������������       �                      @        ������������������������       �                      @        w       |                    @և���X�?             @       x       {                 �UA@���Q��?             @       y       z                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ~       �                     �?�����?:            �V@              �                    �?����X�?5             U@       �       �                    �?=QcG��?            �G@       ������������������������       �                    �B@        �       �                 Ъ�c@�z�G��?             $@       �       �                   �>@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    @��J�fj�?            �B@       �       �                    �?X�<ݚ�?             B@       �       �                    �?X�Cc�?             <@       �       �                    �?8�A�0��?             6@       �       �                   �7@��
ц��?             *@        ������������������������       �                      @        �       �                   �;@�eP*L��?             &@        ������������������������       �                     @        �       �                 p�w@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�q�q�?             "@       �       �                 03�U@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?r�q��?             @       �       �                 �̾w@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 �̰f@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        �       �                    @
�[%G�?�            x@        �       �                    �?���@M^�?             ?@        ������������������������       �                     @        �       �                 @3�4@      �?             8@        ������������������������       �                     &@        �       �                    �?$�q-�?             *@        ������������������������       �                     @        �       �                 ��A>@�����H�?             "@        ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                      @        �       �                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ���@�������?�             v@        �       �                   �=@����-T�?R             _@       �       �                   �<@v�C��?@            �X@       �       �                    �?�q�Q�??             X@        �       �                    �?D�n�3�?             3@        ������������������������       �                     @        �       �                    9@և���X�?	             ,@        �       �                   �1@      �?              @        ������������������������       �                     �?        �       �                 ��y@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                 ���@r�q��?             @        ������������������������       �                      @        �       �                   @<@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        �       �                    �?�w�r��?3            @S@        �       �                    �?      �?             8@       �       �                   �3@��<b���?             7@        �       �                 �?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    8@R���Q�?             4@        ������������������������       �                     @        �       �                   �:@�θ�?             *@        ������������������������       �                      @        �       �                  ��@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     �?        �       �                    �?f1r��g�?#            �J@       �       �                 ��@X�EQ]N�?            �E@        �       �                    6@      �?              @        ������������������������       �                     @        �       �                   �;@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �? >�֕�?            �A@        ������������������������       �                     &@        �       �                    :@�8��8��?             8@       ������������������������       �                     3@        �       �                  s@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                 �&B@�z�G��?             $@        �       �                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �@@`2U0*��?             9@        �       �                   �?@z�G�z�?             @        ������������������������       �                     @        �       �                 �Y5@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     4@        �       �                    �?��t��?�            �l@        �       �                 �?�-@����>�?            �B@        ������������������������       �                     .@        �       �                 03�7@�eP*L��?             6@       �       �                    �?j���� �?             1@       �       �                  �v6@���|���?             &@       �       �                    �?�z�G��?             $@        ������������������������       �                     @        �       �                  �2@      �?             @       �       �                    �?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       4                   @ː����?y             h@       �                       0S�&@�t����?u            `g@       �                          @t��ճC�?O            �`@       �                         �L@�-�[�?N            ``@       �                          �0@����?M            @`@        ������������������������       �      �?              @                                 �?     �?K             `@                                �?���N8�?J            �_@                                �9@d}h���?             ,@        ������������������������       �                     @                              @3�@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @                              ��Y @������?>             \@       	                        @C@p�|�i�?.             S@       
                         ?@     ��?(             P@       ������������������������       �        !            �H@                              @3�@��S�ۿ?             .@       ������������������������       �                     &@                                �@@      �?             @        ������������������������       �                     �?        ������������������������       �                     @                              @3�@r�q��?             (@                                E@      �?              @                               �C@؇���X�?             @       ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     B@        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?              3                   �?x��}�?&            �K@             &                   �?v�X��?             F@             !                   �?�LQ�1	�?             7@                                  5@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        "      #                �T)D@��S�ۿ?
             .@       ������������������������       �                     (@        $      %                   >@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        '      2                ���4@���N8�?             5@       (      -                   0@      �?             $@        )      *                   �?      �?             @        ������������������������       �                     �?        +      ,                ��L.@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        .      /                03;4@�q�q�?             @        ������������������������       �                     @        0      1                  �7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �        	             &@        ������������������������       �                     @        �t�bh�h*h-K ��h/��R�(KM5KK��h]�BP        |@     �p@     `c@     �e@      8@      @      &@              *@      @      &@      @      $@      @      @      @               @      @      �?      �?      �?      �?                      �?      @              @              �?               @       @               @       @             ``@     �d@      Z@     �Y@     �X@     @V@      @      J@      @      E@      @      @      @      �?      @                      �?              @       @     �A@       @      "@              @       @      @      �?      @      �?      �?              @      �?                      :@              $@     �W@     �B@              @     �W@      @@     �E@      8@     �C@      7@      ?@      6@      @      @       @      @      �?              �?      @              @      �?              @              :@      2@      0@      2@              @      0@      (@      (@      @       @              $@      @              �?      $@      @       @               @      @              @       @              @       @              @      @      @      @       @      @                       @               @      $@               @      �?              �?       @              @      �?      @                      �?     �I@       @      :@      @      @      �?      @      �?       @               @      �?              �?       @              �?              5@      @      .@      @      �?              ,@      @      $@              @      @               @      @      @      @      �?      �?              @      �?       @      �?      �?                       @      @              9@       @      @              2@       @      $@       @       @       @       @                       @       @               @              @      ,@               @      @      @       @       @               @       @              @      @      @       @      �?       @               @      �?               @                       @      ;@      P@      8@      N@      @      F@             �B@      @      @      @       @      @                       @              @      5@      0@      4@      0@      2@      $@      *@      "@      @      @       @              @      @              @      @       @      @                       @      @      @      @      �?      @                      �?               @      @      �?      @      �?      @                      �?      �?               @      @              @       @              �?              @      @      @                      @     Pr@      W@      (@      3@              @      (@      (@              &@      (@      �?      @               @      �?      @              @      �?       @              �?      �?              �?      �?             �q@     @R@     �T@     �D@     �M@      D@     �M@     �B@       @      &@              @       @      @      @      @      �?               @      @       @                      @      @      �?       @              @      �?       @      �?      �?             �I@      :@      @      2@      @      2@       @      �?              �?       @              @      1@              @      @      $@       @              �?      $@      �?                      $@      �?             �F@       @      C@      @      @      @      @               @      @              @       @             �@@       @      &@              6@       @      3@              @       @      @                       @      @      @       @      @       @                      @      @                      @      8@      �?      @      �?      @              �?      �?      �?                      �?      4@             �h@      @@      ;@      $@      .@              (@      $@      @      $@      @      @      @      @      @              @      @       @      @              @       @              �?                      �?              @      @             `e@      6@     �d@      6@     �^@      "@     �^@       @     �^@      @      �?      �?     �^@      @      ^@      @      &@      @      @              @      @              @      @             @[@      @     @R@      @     �O@      �?     �H@              ,@      �?      &@              @      �?              �?      @              $@       @      @       @      @      �?      @      �?      @                      �?      @              B@               @                      �?              �?      E@      *@      ?@      *@      .@       @      �?      @      �?                      @      ,@      �?      (@               @      �?       @                      �?      0@      @      @      @      �?      @              �?      �?       @      �?                       @      @       @      @              �?       @      �?                       @      &@              &@              @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ5�;5hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B@E         �                    �?@cF �?�           @�@              	                    /@R�E"��?_           8�@                                   �?���!pc�?             &@                               �y.@z�G�z�?             $@       ������������������������       �                     @                                   )@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        
       G                    �?j[Ԓe�?Y           ��@                                   �?RE��A�?[            �b@                                    @ i���t�?            �H@        ������������������������       �                     :@                                  �5@��<b���?             7@        ������������������������       �                     @                                   �?ףp=
�?             4@                                  �?      �?
             0@        ������������������������       �                     @                                   9@8�Z$���?             *@        ������������������������       �                     �?                                ���@r�q��?             (@        ������������������������       �                     �?                                ���@�C��2(�?             &@        ������������������������       �                     @                                �&B@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     @               :                    �?��x_F-�?<            �Y@              1                    �?�Q��k�?.             T@              *                 ��>@@�0�!��?            �I@               )                  A7@��-�=��?            �C@       !       (                 83�0@      �?             @@       "       #                   �6@��a�n`�?             ?@        ������������������������       �                      @        $       %                   �<@XB���?             =@       ������������������������       �                     4@        &       '                   �=@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        +       0                   �A@�q�q�?             (@       ,       /                    >@      �?              @       -       .                 ���Z@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        2       3                  ��@\-��p�?             =@        ������������������������       �                     $@        4       9                    >@���y4F�?             3@       5       8                   �<@������?             .@       6       7                 ��(@d}h���?             ,@       ������������������������       ��z�G��?             $@        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ;       F                    �?�X����?             6@       <       =                 ��`E@b�2�tk�?             2@        ������������������������       �                     "@        >       ?                   �5@�<ݚ�?             "@        ������������������������       �                     �?        @       A                   �:@      �?              @        ������������������������       �                     @        B       E                 ��hU@      �?             @       C       D                    C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        H       �                 03�S@�*I�?�            Px@       I       n                    �?�`��ie�?�            �v@        J       a                   �:@(���X�?,            @Q@        K       L                 pf�@�P�*�?             ?@        ������������������������       �                      @        M       `                    �?\X��t�?             7@       N       [                    �?�eP*L��?             6@       O       P                     @և���X�?             ,@        ������������������������       �                     @        Q       Z                   �6@���!pc�?             &@       R       U                    3@      �?              @        S       T                 ��!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        V       W                    5@�q�q�?             @        ������������������������       �                     �?        X       Y                 �̜!@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        \       ]                 �̬)@      �?              @       ������������������������       �                     @        ^       _                 @3�/@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        b       m                   @G@>A�F<�?             C@       c       l                 `f�&@�������?             >@        d       e                   �;@�<ݚ�?             "@        ������������������������       �                     �?        f       k                    �?      �?              @       g       h                 `�X!@r�q��?             @       ������������������������       �                     @        i       j                  SE"@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     5@        ������������������������       �                      @        o       �                     �?l������?�            �r@        p       s                 03k:@��s����?             E@        q       r                   �9@      �?             @       ������������������������       �                     @        ������������������������       �                     @        t       �                    �?4?,R��?             B@       u       �                   �<@     ��?             @@        v       w                   �;@      �?	             $@        ������������������������       �                     �?        x                        ��yC@X�<ݚ�?             "@       y       z                 `fF<@և���X�?             @        ������������������������       ��q�q�?             @        {       |                   �>@      �?             @        ������������������������       �                      @        }       ~                   �@@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     6@        ������������������������       �                     @        �       �                     @      �?�             p@        �       �                   �@@��?^�k�?-            �Q@       ������������������������       �                     D@        �       �                   @A@��S�ۿ?             >@        ������������������������       �      �?              @        �       �                   �E@h�����?             <@        �       �                   �3@$�q-�?             *@       �       �                   �'@      �?              @        ������������������������       �                     @        �       �                   @D@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �        
             .@        �       �                 �T)D@㺦���?x            @g@       �       �                   �0@�D����?u            �f@        �       �                 pf�@�q�q�?             @        ������������������������       �                     �?        �       �                 pFD!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �<@8�be��?r            @f@       �       �                  ��	@     8�?O             `@        �       �                    6@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �? ;=֦��?M            �^@       �       �                   �:@��9J���?B             Z@       �       �                 �1@P����?&            �M@        �       �                 �?$@���7�?             6@       ������������������������       �                     3@        �       �                   �5@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                    �B@        �       �                   �;@`Ӹ����?            �F@        ������������������������       �                     �?        �       �                 �?$@`���i��?             F@        �       �                 pf�@ףp=
�?             $@       ������������������������       �                      @        ������������������������       �      �?              @        ������������������������       �                     A@        ������������������������       �                     2@        �       �                    �?H%u��?#             I@       �       �                   @@@      �?!             H@        �       �                   �>@�q�q�?             (@        �       �                   �=@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �?�@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                 �?�@������?             B@       ������������������������       �                     3@        �       �                   �E@�IєX�?             1@       ������������������������       �                     *@        �       �                   �F@      �?             @        �       �                 @3�@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    ;@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�C��2(�?             6@       ������������������������       �                     4@        ������������������������       �                      @        �       �                     @�4��'��?k             d@        �       �                    �?x�(�3��?2            @S@       �       �                   �2@�q�q�?/            @Q@        �       �                    @P���Q�?             4@        �       �                    �?؇���X�?             @       ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     *@        �       �                    �?Tt�ó��?!            �H@       �       �                    �? �Cc}�?             <@       ������������������������       �        
             2@        �       �                    �?�z�G��?             $@        ������������������������       �                     �?        �       �                   �8@�q�q�?             "@        ������������������������       �                     @        �       �                     �?      �?             @       �       �                   �>@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?�����?             5@        ������������������������       �                      @        �       �                    �?8�Z$���?
             *@       ������������������������       �                     "@        �       �                    �?      �?             @        ������������������������       �                     �?        �       �                     �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �                          �?�q�q�?9             U@       �       �                    @X�<ݚ�?            �F@        �       �                 P��%@"pc�
�?             &@        ������������������������       �                     �?        �       �                 0C�7@ףp=
�?             $@       ������������������������       �                      @        �       �                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�!���?             A@        �       �                    @r�q��?             @       �       �                   �<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �                       ���4@d}h���?             <@        �                           @���Q��?             $@       �       �                    �?X�<ݚ�?             "@       �       �                    >@      �?             @       �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     2@                                 �?x�����?            �C@                              =
�@      �?             @        ������������������������       �                      @                              ��&@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        	      
                   �?؇���X�?            �A@        ������������������������       �                     @                                  @r�q��?             >@                                 �?������?	             .@        ������������������������       �                     @                                 &@���|���?             &@        ������������������������       �                     @        ������������������������       �                     @                                 @��S�ۿ?
             .@                              ���A@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     *@        �t�b�`)     h�h*h-K ��h/��R�(KMKK��h]�BP       }@     �n@      x@     �d@      @       @       @       @              @       @       @       @                       @      �?             �w@     �c@     �U@      P@      @      F@              :@      @      2@      @               @      2@       @      ,@              @       @      &@              �?       @      $@      �?              �?      $@              @      �?      @      �?       @              �?              @     �T@      4@     �P@      *@      E@      "@     �A@      @      <@      @      <@      @               @      <@      �?      4@               @      �?              �?       @                      �?      @              @      @      @      @      @      �?              �?      @                      @      @              9@      @      $@              .@      @      &@      @      &@      @      @      @      @                      �?      @              .@      @      &@      @      "@               @      @      �?              �?      @              @      �?      @      �?      �?      �?                      �?               @      @             �r@     @W@     `r@     @R@      4@     �H@      *@      2@               @      *@      $@      (@      $@       @      @              @       @      @      @      @      �?      �?      �?                      �?      @       @      �?              @       @               @      @              @              @      @      @              �?      @              @      �?              �?              @      ?@      @      7@      @       @              �?      @      �?      @      �?      @              �?      �?              �?      �?               @                      5@               @      q@      8@      A@       @      @      @      @                      @      ?@      @      ;@      @      @      @              �?      @      @      @      @       @      �?      �?      @               @      �?      �?      �?                      �?       @              6@              @              n@      0@      Q@       @      D@              <@       @      �?      �?      ;@      �?      (@      �?      @      �?      @              @      �?      �?               @      �?      @              .@             �e@      ,@      e@      (@       @      �?      �?              �?      �?              �?      �?             �d@      &@     �^@      @      @       @      @                       @     �]@      @     @Y@      @      M@      �?      5@      �?      3@               @      �?              �?       @             �B@             �E@       @              �?     �E@      �?      "@      �?       @              �?      �?      A@              2@              F@      @      E@      @      @      @      @      �?              �?      @               @      @       @                      @     �A@      �?      3@              0@      �?      *@              @      �?      �?      �?              �?      �?               @               @              @       @               @      @               @      4@              4@       @             �S@     �T@      7@      K@      7@      G@      �?      3@      �?      @              @      �?       @      �?                       @              *@      6@      ;@      @      9@              2@      @      @              �?      @      @              @      @      @      @       @      @                       @              �?      3@       @       @              &@       @      "@               @       @      �?              �?       @               @      �?                       @      L@      <@      9@      4@       @      "@      �?              �?      "@               @      �?      �?      �?                      �?      7@      &@      �?      @      �?       @      �?                       @              @      6@      @      @      @      @      @      �?      @      �?      �?              �?      �?                       @      @       @      @                       @              �?      2@              ?@       @      �?      @               @      �?      �?      �?                      �?      >@      @      @              9@      @      &@      @      @              @      @              @      @              ,@      �?      �?      �?              �?      �?              *@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJi4�hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM_huh*h-K ��h/��R�(KM_��h|�B�W         �                     @�)�>_M�?�           @�@               s                    �?0�矆��?�            �t@              h                   �I@r�q��?�             h@              /                     �?j4�����?r             e@               *                    �?"+q��?4            @S@                                 �;@և���X�?,            �O@        ������������������������       �                      @                                  �=@D7�J��?&            �K@        	                        `ffP@�q�q�?             5@       
                          �<@�z�G��?             4@                                  �?�q�q�?             2@                                �ܵ<@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?                                  �>@�q�q�?             .@                               `fF<@X�<ݚ�?             "@                               �̌*@z�G�z�?             @        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?                                   �?h+�v:�?             A@                                   G@�IєX�?             1@       ������������������������       �        
             0@        ������������������������       �                     �?               #                 `f&;@�t����?             1@                                ��I*@      �?              @        ������������������������       �                     @                                    D@z�G�z�?             @        ������������������������       �                     @        !       "                    H@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        $       )                    �?�����H�?             "@       %       &                    =@r�q��?             @        ������������������������       �                     @        '       (                   �A@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        +       ,                    �?����X�?             ,@        ������������������������       �                     @        -       .                 @��v@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        0       5                    �?��c:�?>             W@        1       2                 `��,@���Q��?             $@        ������������������������       �                     @        3       4                    �?�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        6       W                   �C@hP�vCu�?8            �T@       7       T                    �?:ɨ��?-            �P@       8       ?                 `fF)@�BbΊ�?'             M@        9       :                    @�����H�?             2@        ������������������������       �                      @        ;       <                   �:@      �?             0@        ������������������������       �                     @        =       >                    �?�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        @       S                   �J@�G�z�?             D@       A       D                   �;@*O���?             B@        B       C                    �?8�Z$���?	             *@        ������������������������       �      �?             @        ������������������������       �                     "@        E       R                   �=@
;&����?             7@       F       Q                   �B@���Q��?             4@       G       H                    �?��.k���?             1@        ������������������������       �                     @        I       L                    =@      �?             (@        J       K                   �*@      �?             @        ������������������������       �                      @        ������������������������       �                      @        M       N                    @@      �?              @        ������������������������       �                     @        O       P                   �3@z�G�z�?             @       ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        U       V                    �?      �?              @       ������������������������       �                     @        ������������������������       �                     @        X       g                   @I@      �?             0@       Y       f                   �6@z�G�z�?
             .@       Z       a                   �,@؇���X�?	             ,@       [       \                   �'@�C��2(�?             &@        ������������������������       �                     @        ]       `                   �*@      �?              @       ^       _                    �?؇���X�?             @        ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                     �?        b       e                    �?�q�q�?             @       c       d                   �.@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        i       r                     �?�㙢�c�?             7@       j       q                 ��{P@������?             1@       k       l                    �?�r����?
             .@        ������������������������       �                      @        m       n                    �?8�Z$���?	             *@        ������������������������       �                     �?        o       p                    R@�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        t       u                    2@�>z���?R             a@        ������������������������       �                     .@        v       �                  ��S@��Fh�?E            @^@       w       x                    �?ؤ�u��?1            �T@       ������������������������       �                     G@        y       �                     �?����>�?            �B@        z       {                  x#J@�n_Y�K�?             *@        ������������������������       �                     @        |       }                    �?      �?              @        ������������������������       �                      @        ~                           7@      �?             @        ������������������������       �                      @        �       �                   �J@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    @@�q�q�?             8@        �       �                   �?@�n_Y�K�?             *@       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        	             &@        �       �                    �?�\��N��?             C@        �       �                    8@�8��8��?             (@        ������������������������       �                     @        �       �                 ���`@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?R�}e�.�?             :@       �       �                   �G@��S���?             .@       �       �                   �:@�z�G��?             $@        ������������������������       �                     �?        �       �                 03�U@�<ݚ�?             "@       ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                 `f^@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        �       R                  @B@�q�q*�?�             x@       �       E                   �?������?�            pu@       �       �                   �0@\N�pV�?�            �r@        �       �                    �?�4�����?             ?@       �       �                    �?�q�q�?             8@        �       �                    �?�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        �       �                   �&@���Q��?	             .@       �       �                 P��@      �?              @        ������������������������       �                      @        �       �                 �̌!@      �?             @        ������������������������       �      �?             @        ������������������������       �                      @        �       �                     @؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 ��\"@և���X�?             @        ������������������������       �                     �?        �       �                    �?�q�q�?             @        �       �                 �&�)@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �                       `�X.@b�28ƿ�?�            �p@       �       �                    �?�����?�            �k@        �       �                 @3�@
;&����?             G@       �       �                    �?�q�q�?            �@@        ������������������������       �                     @        �       �                    �?����"�?             =@        �       �                    9@      �?	             0@        ������������������������       �                     �?        �       �                  ��@���Q��?             .@        ������������������������       �                     @        �       �                 �&B@"pc�
�?             &@       �       �                 ���@�<ݚ�?             "@        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                      @        �       �                    �?�n_Y�K�?	             *@       �       �                   �9@�q�q�?             (@       �       �                   �6@և���X�?             @        ������������������������       �                      @        �       �                 pf�@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?8�Z$���?
             *@       �       �                    =@�8��8��?	             (@       ������������������������       �                     &@        ������������������������       �                     �?        ������������������������       �                     �?        �                         �<@ �<#�?o            �e@       �       �                 �1@�#-���?V            �a@        �       �                 �?$@R���Q�?$             N@       �       �                   �3@      �?!             L@        ������������������������       �                     (@        �       �                 �Y�@fP*L��?             F@        �       �                    5@���N8�?             5@        �       �                 �{@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?r�q��?             2@       �       �                    �?�r����?	             .@       �       �                 ���@r�q��?             (@        ������������������������       �                     @        ������������������������       �����X�?             @        ������������������������       �                     @        �       �                 ���@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?���}<S�?             7@        �       �                   �:@�C��2(�?             &@        ������������������������       �                     �?        �       �                 03�@ףp=
�?             $@        ������������������������       �                     �?        �       �                    �?�����H�?             "@       ������������������������       �r�q��?             @        ������������������������       �                     @        �       �                 ��@�8��8��?             (@       ������������������������       �                     $@        �       �                    ;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �;@      �?             @       ������������������������       �                      @        ������������������������       �                      @        �       �                   �4@x�G�z�?2             T@        �       �                   �3@�����H�?
             2@        ������������������������       �                     (@        �       �                 @3�@�q�q�?             @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                 ��) @0�z��?�?(             O@       ������������������������       �                     G@        �                           �?      �?             0@       �       �                 pf� @@4և���?
             ,@        ������������������������       �                     �?        ������������������������       �        	             *@        ������������������������       �                      @                                 @����X�?            �A@        ������������������������       �                     @                                 �?J�8���?             =@                                 ?@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @                              @3�@���!pc�?             6@        	      
                  �?@���Q��?             $@        ������������������������       �                      @                                �@      �?              @        ������������������������       �                     �?                                @@@և���X�?             @                             �?�@      �?             @        ������������������������       �                     �?        ������������������������       ����Q��?             @        ������������������������       �                     �?                                �=@r�q��?	             (@                              �̌!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                @@@ףp=
�?             $@                                 ?@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @                                 3@      �?!             I@        ������������������������       �                     @              (                   �?JJ����?             �G@              '                   �?�����H�?             "@             &                   �?      �?              @              %                   @z�G�z�?             @       !      $                  �<@�q�q�?             @       "      #                 S�2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        )      D                   A@�s��:��?             C@       *      3                   �?���Q��?            �A@        +      2                ���5@����X�?	             ,@       ,      -                   �?�C��2(�?             &@        ������������������������       �                     @        .      /                ��Y1@      �?              @       ������������������������       �                     @        0      1                03C3@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        4      A                   ?@��s����?             5@       5      8                   ;@      �?             0@        6      7                   �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        9      @                  @<@�8��8��?             (@       :      ;                   �?�����H�?             "@        ������������������������       �                      @        <      ?                   �?؇���X�?             @       =      >                �T�C@r�q��?             @        ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     @        B      C                �TAC@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        F      I                   �?��p\�?            �D@        G      H                   @z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        J      K                   �?�X�<ݺ?             B@        ������������������������       �                     �?        L      Q                   �?��?^�k�?            �A@        M      N                  �0@@4և���?	             ,@       ������������������������       �                     $@        O      P                8#�0@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             5@        S      \                  �N@������?            �D@       T      [                  @F@P�Lt�<�?             C@       U      V                   �?�X�<ݺ?             2@        ������������������������       �                      @        W      X                �?�@      �?             0@        ������������������������       �                     @        Y      Z                  �E@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     4@        ]      ^                ��\!@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �t�bh�h*h-K ��h/��R�(KM_KK��h]�B�       `{@      q@     �b@      f@      Z@      V@     @U@      U@      ?@      G@      ;@      B@               @      ;@      <@      ,@      @      ,@      @      (@      @       @      �?       @                      �?      $@      @      @      @      @      �?      @              �?      �?              @      @               @                      �?      *@      5@      �?      0@              0@      �?              (@      @      @      @      @              �?      @              @      �?      �?      �?                      �?       @      �?      @      �?      @               @      �?              �?       @              @              @      $@              @      @      @      @                      @      K@      C@      @      @              @      @       @      @                       @      I@      @@      G@      4@     �E@      .@      0@       @       @              ,@       @      @              @       @               @      @              ;@      *@      7@      *@      &@       @       @       @      "@              (@      &@      (@       @      "@       @              @      "@      @       @       @               @       @              @      �?      @              @      �?       @      �?       @              @                      @      @              @      @              @      @              @      (@      @      (@       @      (@      �?      $@              @      �?      @      �?      @              @      �?       @              �?      �?       @      �?      �?      �?                      �?              �?      �?              �?              3@      @      *@      @      *@       @       @              &@       @              �?      &@      �?      &@                      �?               @      @             �G@     @V@              .@     �G@     �R@      ;@      L@              G@      ;@      $@       @      @      @              @      @               @      @      @       @              �?      @              @      �?              3@      @       @      @       @                      @      &@              4@      2@      �?      &@              @      �?      @              @      �?              3@      @       @      @      @      @              �?      @       @      @               @       @               @       @              �?      @      �?                      @      &@             �q@     @X@      o@     �W@     @j@      W@      $@      5@      @      1@      �?       @               @      �?              @      "@      @      @       @              @      @      �?      @       @              �?      @              @      �?              @      @      �?               @      @       @       @               @       @                       @      i@     �Q@     �e@      G@      6@      8@      &@      6@              @      &@      2@      @      $@              �?      @      "@      @               @      "@       @      @              �?       @      @               @      @       @      @       @      @      @               @      @      �?              �?      @                      @      �?              &@       @      &@      �?      &@                      �?              �?      c@      6@      `@      (@     �I@      "@     �H@      @      (@             �B@      @      0@      @      �?       @      �?                       @      .@      @      *@       @      $@       @      @              @       @      @               @      �?       @                      �?      5@       @      $@      �?      �?              "@      �?      �?               @      �?      @      �?      @              &@      �?      $@              �?      �?      �?                      �?       @       @               @       @             @S@      @      0@       @      (@              @       @      �?       @      �?                       @      @             �N@      �?      G@              .@      �?      *@      �?              �?      *@               @              9@      $@      @              3@      $@      @      @              @      @              0@      @      @      @       @              @      @              �?      @      @      @      @      �?               @      @      �?              $@       @      �?      �?      �?                      �?      "@      �?      @      �?      @                      �?      @              9@      9@      @              6@      9@      �?       @      �?      @      �?      @      �?       @      �?      �?      �?                      �?              �?               @              @              �?      5@      1@      5@      ,@      @      $@      �?      $@              @      �?      @              @      �?      @      �?                      @      @              1@      @      ,@       @      @      �?              �?      @              &@      �?       @      �?       @              @      �?      @      �?      @               @      �?      �?              @              @       @      @                       @              @      C@      @      @      �?      @                      �?      A@       @              �?      A@      �?      *@      �?      $@              @      �?              �?      @              5@             �C@       @     �B@      �?      1@      �?       @              .@      �?      @               @      �?       @                      �?      4@               @      �?       @                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�ThG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM-huh*h-K ��h/��R�(KM-��h|�B@K         x                     @z����?�           @�@                                   �?�l5wA��?�            ps@                                   �?���?W            �`@              	                   �*@���#�İ?L            �]@                                ��Y)@��2(&�?             6@        ������������������������       �                     @                                   :@     ��?             0@        ������������������������       ����Q��?             @        ������������������������       �                     &@        
                        ���@@�q�q�?A             X@                                  �H@г�wY;�?             A@       ������������������������       �                     :@                                    �?      �?              @                                   K@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        -             O@                                    �?������?             1@                                   �?և���X�?             @        ������������������������       �                     �?                                   *@�q�q�?             @        ������������������������       �                      @                                    @      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     $@                                   (@�7�A�?p             f@        ������������������������       �                     @               1                    �?;���?j             e@               "                 pVAH@     ��?             @@                !                 ���,@�r����?	             .@        ������������������������       �                      @        ������������������������       �                     *@        #       ,                 �U�X@��.k���?             1@       $       %                    �?�<ݚ�?             "@        ������������������������       �                     �?        &       +                    C@      �?              @        '       (                 ��3Q@�q�q�?             @        ������������������������       �                     �?        )       *                   �:@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        -       0                 �̾w@      �?              @       .       /                   �1@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        2       Q                   �@@|���~�?T             a@       3       >                 `fF:@�KM�]�?+             S@       4       5                     �?`'�J�?            �I@        ������������������������       �                     @        6       =                    &@���7�?             F@        7       8                    @�t����?	             1@        ������������������������       �                     @        9       <                   �5@z�G�z�?             $@        :       ;                   �1@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     ;@        ?       @                 `fF<@�+e�X�?             9@        ������������������������       �                      @        A       P                    �?�㙢�c�?             7@       B       C                   @>@�<ݚ�?             2@        ������������������������       �                      @        D       E                   �9@      �?
             0@        ������������������������       �                     @        F       M                    �?�q�q�?             (@       G       H                   `@@�<ݚ�?             "@        ������������������������       �                     �?        I       L                 ��yC@      �?              @        J       K                   �A@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        N       O                   �=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        R       S                    �?��6}��?)            �N@        ������������������������       �                     @        T       m                     �?��h!��?'            �L@       U       V                   �B@��>4և�?             <@        ������������������������       �                     @        W       f                   �J@`�Q��?             9@       X       a                 �T!@@     ��?             0@       Y       `                    H@���Q��?             $@       Z       _                 `f�;@�q�q�?             @       [       \                   @D@      �?             @        ������������������������       �                     �?        ]       ^                 03k:@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     @        b       c                 XfZX@r�q��?             @        ������������������������       �                     @        d       e                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        g       l                    �?�����H�?             "@       h       i                 `fF<@r�q��?             @        ������������������������       �                     @        j       k                   @>@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        n       w                   �*@д>��C�?             =@       o       v                    G@�E��ӭ�?
             2@       p       u                   @D@�q�q�?             (@       q       r                   �'@�<ݚ�?             "@        ������������������������       �                     @        s       t                   @B@�q�q�?             @       ������������������������       ����Q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        	             &@        y       �                    �?1`�N�?�            y@        z       �                   @B@��%��?G            �[@       {       �                    @@x��#���?@             Y@       |       �                    @��C����?>            �W@       }       ~                    @LMc����?4            @T@        ������������������������       �                     @               �                 ��@�EH,���?1            �R@        �       �                    �?�<ݚ�?             2@        ������������������������       �                     @        �       �                   �5@����X�?             ,@        �       �                 ���@���Q��?             @        ������������������������       �                      @        �       �                    �?�q�q�?             @       �       �                  s�@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �9@�����H�?             "@        ������������������������       �                     @        �       �                 ���@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?D�n�3�?"            �L@       �       �                    �?����"�?             =@        �       �                    �?      �?              @       �       �                 `�@1@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �=@����X�?             5@       �       �                    0@      �?             4@        ������������������������       �                     @        �       �                    3@�t����?             1@        �       �                    �?      �?             @       �       �                 ��!@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 pf� @"pc�
�?             &@        �       �                 �?�@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                 �y7+@      �?              @       ������������������������       �                     @        �       �                   �:@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �6@���>4��?             <@        ������������������������       �                     @        �       �                    �?\X��t�?             7@       �       �                    �?����X�?	             ,@       �       �                 ��1@�q�q�?             (@       �       �                    ;@z�G�z�?             $@        �       �                   �8@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                    >@�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        �       �                   -@؇���X�?
             ,@        ������������������������       �                     �?        �       �                    �?$�q-�?	             *@        ������������������������       �                     @        �       �                 ��T?@؇���X�?             @        ������������������������       �                     @        �       �                    %@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     &@        �       �                    '@Riv����?�             r@        �       �                     @և���X�?
             5@        ������������������������       �                     &@        �       �                    �?ףp=
�?             $@        ������������������������       �                     @        �       �                     @      �?             @        ������������������������       �                      @        �       �                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �                       ���5@Pz�
r��?�            �p@       �       �                   �	@���I�?�            @n@        �       �                    6@�q�q�?             @        ������������������������       �                     �?        �       �                   �>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �                          �?`.��A��?�            �m@       �                          �?��ϭ�*�?�             m@       �       �                   �:@���d���?~            `i@        �       �                 03�@0�,���?*            �P@        �       �                 �̌@؇���X�?             @       ������������������������       �                     @        �       �                   �7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �0@ �.�?Ƞ?%             N@        �       �                 pFD!@      �?              @       �       �                 pf�@z�G�z�?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                      J@        �       �                  s�@���� �?T             a@        �       �                    �?P�Lt�<�?             C@       ������������������������       �                     9@        �       �                 033@$�q-�?             *@        �       �                   �>@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   �@؇���X�?<            �X@        �       �                 ��@�q�q�?             8@       �       �                    >@������?	             1@       �       �                   �<@�q�q�?             (@       ������������������������       �z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                     @        �       �                    D@և���X�?             @       �       �                   �=@z�G�z�?             @        ������������������������       �                      @        �       �                 �&B@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �                          �?�L���?.            �R@       �       �                   �;@@�j;��?,            �Q@        ������������������������       �                      @        �       �                 �?�@p��%���?+            @Q@        ������������������������       �                     8@        �                         @B@�:�^���?            �F@                                @<@ >�֕�?            �A@                             ��) @�����?             5@       ������������������������       �                     .@                              pf� @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        
             ,@                                @D@z�G�z�?             $@        ������������������������       �                     �?        	      
                @3�@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                 �?ܷ��?��?             =@                                �?P���Q�?             4@        ������������������������       �                     @                                �8@��S�ۿ?	             .@        ������������������������       �                      @                              �&B@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @                                 7@�<ݚ�?             "@                             茘'@���Q��?             @        ������������������������       �                      @                                 2@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @                                  �?X�<ݚ�?             ;@                                 �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        !      "                   9@�q�q�?             5@        ������������������������       �                     @        #      ,                p�O@b�2�tk�?	             2@       $      +                   �?��
ц��?             *@       %      &                �T)D@���|���?             &@        ������������������������       �                     �?        '      *                   >@�z�G��?             $@       (      )                   ;@և���X�?             @        ������������������������       �                     �?        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �t�bh�h*h-K ��h/��R�(KM-KK��h]�B�       �{@     �p@     �a@      e@       @     �_@      @     �\@      @      3@              @      @      *@      @       @              &@      �?     �W@      �?     �@@              :@      �?      @      �?      @      �?                      @              @              O@      @      *@      @      @              �?      @       @       @               @       @       @                       @              $@     �`@      E@              @     �`@     �A@      5@      &@      *@       @               @      *@               @      "@       @      @      �?              �?      @      �?       @              �?      �?      �?              �?      �?                      @      @       @      @      �?              �?      @                      �?     @\@      8@      Q@       @     �H@       @      @              E@       @      .@       @      @               @       @       @       @       @                       @      @              ;@              3@      @               @      3@      @      ,@      @       @              (@      @      @               @      @      @       @              �?      @      �?       @      �?       @                      �?      @              �?       @               @      �?              @             �F@      0@      @             �D@      0@      1@      &@              @      1@       @      "@      @      @      @      @       @       @       @      �?              �?       @              �?      �?      �?       @                      @      @      �?      @              �?      �?              �?      �?               @      �?      @      �?      @               @      �?              �?       @              @              8@      @      *@      @      @      @      @       @      @              @       @      @       @      �?                      @      @              &@             s@      X@      N@     �I@     �H@     �I@     �H@      G@     �B@      F@              @     �B@      C@      @      ,@              @      @      $@      @       @       @              �?       @      �?      �?              �?      �?                      �?      �?       @              @      �?      @      �?                      @     �@@      8@      2@      &@      @      @      @       @      @                       @              @      .@      @      .@      @      @              (@      @      @      @      @      �?      @                      �?               @      "@       @       @      �?       @                      �?      @      �?      @               @      �?              �?       @                      �?      .@      *@      @              $@      *@      @      $@      @       @       @       @       @       @               @       @                      @       @                       @      @      @      @                      @      (@       @              �?      (@      �?      @              @      �?      @              @      �?              �?      @                      @      &@             �n@     �F@      "@      (@              &@      "@      �?      @              @      �?       @              �?      �?              �?      �?             �m@     �@@     �k@      5@       @      �?      �?              �?      �?              �?      �?             `k@      4@     �j@      4@     @g@      1@     @P@       @      @      �?      @               @      �?              �?       @             �M@      �?      @      �?      @      �?       @               @      �?      @              J@             @^@      .@     �B@      �?      9@              (@      �?      @      �?              �?      @               @              U@      ,@      0@       @      *@      @       @      @       @       @               @      @              @      @      �?      @               @      �?       @      �?                       @       @              Q@      @     @P@      @               @     @P@      @      8@             �D@      @     �@@       @      3@       @      .@              @       @               @      @              ,@               @       @              �?       @      �?              �?       @              @              :@      @      3@      �?      @              ,@      �?       @              @      �?              �?      @              @       @      @       @       @              �?       @      �?                       @      @              @              .@      (@      �?      @      �?                      @      ,@      @      @              &@      @      @      @      @      @      �?              @      @      @      @              �?      @      @              @       @              @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ5�R/hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM#huh*h-K ��h/��R�(KM#��h|�B�H         R                    �?4�<����?�           @�@                                    @d�� z�?�            `n@                                  �?P�� �?Q            @`@                                  �?��FM ò?C            @Z@               
                    �?      �?             @@              	                 hލC@ףp=
�?             4@                                `v7<@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        	             *@        ������������������������       �                     (@                                   6@��pBI�?0            @R@                                   �?�C��2(�?             6@        ������������������������       �                     @                                   �?�KM�]�?             3@                                 �;@�t����?             1@                                   1@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     (@        ������������������������       �                      @        ������������������������       �        #            �I@                                ���`@z�G�z�?             9@       ������������������������       �        
             1@                                   �?      �?              @        ������������������������       �                     @        ������������������������       �                     @               Q                 �A7@+Y���?G            @\@              B                    .@<SvLB�?9             W@              )                 ��@�'�=z��?(            �P@               (                    �?      �?             4@               !                    9@r�q��?             2@        ������������������������       �                     @        "       %                  ��@���!pc�?             &@        #       $                 0��@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        &       '                 ���@      �?              @        ������������������������       �                     @        ������������������������       �z�G�z�?             @        ������������������������       �                      @        *       +                    �?nM`����?             G@        ������������������������       �                     @        ,       -                 0�w@H�z�G�?             D@        ������������������������       �                     @        .       A                    �?      �?             A@       /       @                    �?*;L]n�?             >@       0       5                 pF @\X��t�?             7@        1       2                    �?      �?              @       ������������������������       �                     @        3       4                 �?�@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        6       ;                    =@���Q��?
             .@       7       :                    �?z�G�z�?             $@       8       9                    3@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        <       =                   �@@z�G�z�?             @        ������������������������       �                      @        >       ?                    I@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        C       N                    @���B���?             :@       D       E                 03�1@�LQ�1	�?             7@        ������������������������       �                      @        F       G                   �<@z�G�z�?
             .@       ������������������������       �                     "@        H       M                   �@@      �?             @       I       J                 03C3@      �?             @        ������������������������       �                      @        K       L                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        O       P                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     5@        S                          �?��%n��?&           P}@       T                         @S@�7�iU�?�            Px@       U       �                     �?ʩ�ժ�?�            0x@        V       i                 ��9L@��W3�?-            �Q@       W       h                    �?������?            �F@       X       [                    ?@�z�G��?             D@        Y       Z                   �;@�����H�?
             2@        ������������������������       �                      @        ������������������������       �        	             0@        \       g                   �B@�eP*L��?             6@       ]       ^                   �9@X�<ݚ�?             2@        ������������������������       �                     �?        _       b                    �?j���� �?             1@        `       a                   �L@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        c       f                    @@և���X�?
             ,@       d       e                    L@�q�q�?             (@       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        j       k                   �7@      �?             :@        ������������������������       �                     @        l       m                   �;@\X��t�?             7@        ������������������������       �                     @        n                           �?X�<ݚ�?             2@       o       p                 03�M@��.k���?             1@        ������������������������       �                     @        q       r                    @@X�Cc�?
             ,@        ������������������������       �                     @        s       t                    �?      �?             $@        ������������������������       �                      @        u       x                 ЈrS@      �?              @        v       w                   �G@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        y       z                    �?z�G�z�?             @        ������������������������       �                     �?        {       |                   �B@      �?             @        ������������������������       �                      @        }       ~                   �D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?l�YS��?�            �s@       �       �                    A@��FA6�?�             s@       �       �                    �? E=��H�?�             o@       �       �                 ��@�������?�            �j@        �       �                   �;@     ��?             0@        �       �                 ���@�<ݚ�?             "@       �       �                 033@�q�q�?             @       �       �                 `f�@z�G�z�?             @       �       �                    6@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 �?�@�q��/��?{            �h@        �       �                   �<@p�eU}�?=            �Y@       �       �                   �5@h�����?3             U@        ������������������������       �        	             1@        �       �                    �?�����?*            �P@        �       �                   �7@��S�ۿ?             >@        �       �                 ���@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �? 7���B�?             ;@       ������������������������       �                     *@        �       �                  s�@@4և���?             ,@        ������������������������       �                     @        �       �                 ��(@�C��2(�?             &@       ������������������������       �ףp=
�?             $@        ������������������������       �                     �?        �       �                    ;@�?�|�?            �B@        ������������������������       �                     &@        �       �                  sW@ ��WV�?             :@        �       �                 pf�@ףp=
�?             $@       ������������������������       �                      @        ������������������������       �      �?              @        ������������������������       �        	             0@        �       �                    �?�S����?
             3@        ������������������������       �                     �?        �       �                    �?�����H�?	             2@        �       �                    >@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �@$�q-�?             *@        �       �                 �&B@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �@@�n`���?>            @W@       �       �                     @��zi��?=            �V@        �       �                   �(@ �q�q�?             8@        ������������������������       �                     $@        �       �                   �*@@4և���?             ,@        �       �                   �:@z�G�z�?             @       ������������������������       �                     @        �       �                    =@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        �       �                    �?��ga�=�?+            �P@        �       �                    ;@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �7@�������?&             N@        �       �                 ��Y @؇���X�?             5@        �       �                   �3@      �?             (@       �       �                   �1@և���X�?             @        ������������������������       �      �?             @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     "@        �       �                 @3�@�(�Tw��?            �C@        ������������������������       �                      @        �       �                 ��) @���"͏�?            �B@        ������������������������       �                     .@        �       �                   �>@8�A�0��?             6@       �       �                 �̜!@     ��?	             0@        ������������������������       �                     @        �       �                    ;@���|���?             &@        ������������������������       �                      @        �       �                   �<@�<ݚ�?             "@       �       �                 �!&B@      �?              @       ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�8��8��?             B@        ������������������������       �                      @        �       �                 ��l#@ �Cc}�?             <@        �       �                 P�@�<ݚ�?             "@       �       �                   �7@      �?              @       ������������������������       �                     @        �       �                 �&B@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �7@�}�+r��?
             3@       ������������������������       �                     ,@        �       �                   �<@z�G�z�?             @        ������������������������       �                      @        �       �                   �@@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �N@�8���?$             M@       �       �                    �?�&=�w��?             �J@       �       �                   @C@ ��WV�?             J@        ������������������������       �        	             4@        �       �                    �?      �?             @@        ������������������������       �                     @        �       �                   �E@ 	��p�?             =@        �       �                     @�<ݚ�?             "@        �       �                   @D@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 �?�@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     4@        ������������������������       �                     �?        �       �                     @z�G�z�?             @        �       �                   �P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �                           ;@z�G�z�?             $@        ������������������������       �                     @                                 �?����X�?             @                                 �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @              "                   @�z�G��?0             T@                                @��cv�?.            @S@        	                         @�ՙ/�?             5@       
                          @X�<ݚ�?
             2@        ������������������������       �                     $@        ������������������������       �                      @        ������������������������       �                     @              !                    @����>4�?#             L@                                6@�%^�?            �E@                                �0@r�q��?             @                                 )@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                 �?�MI8d�?            �B@        ������������������������       �                     (@                                   �?�+e�X�?             9@                               x�N@      �?             (@        ������������������������       �                      @                               D�\@���Q��?             $@                             `f�R@      �?              @        ������������������������       �                     @                              03�S@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     *@        ������������������������       �                     *@        ������������������������       �                     @        �t�b��r      h�h*h-K ��h/��R�(KM#KK��h]�B0        |@     �p@     @Q@     �e@      "@     @^@      @     @Y@       @      >@       @      2@       @      @              @       @                      *@              (@       @     �Q@       @      4@              @       @      1@       @      .@       @      @              @       @                      (@               @             �I@      @      4@              1@      @      @      @                      @      N@     �J@     �C@     �J@      A@      @@      @      .@      @      .@              @      @       @       @      �?              �?       @              �?      @              @      �?      @       @              =@      1@      @              7@      1@      @              1@      1@      1@      *@      $@      *@      �?      @              @      �?      �?      �?                      �?      "@      @       @       @       @      �?              �?       @                      �?      �?      @               @      �?       @      �?                       @      @                      @      @      5@      @      4@               @      @      (@              "@      @      @      @      �?       @              �?      �?              �?      �?                       @       @      �?              �?       @              5@             �w@     �V@     0t@     �P@     0t@      P@      G@      9@     �@@      (@      <@      (@      0@       @               @      0@              (@      $@       @      $@      �?              @      $@      �?       @               @      �?              @       @      @       @               @      @               @              @              @              *@      *@      @              $@      *@              @      $@       @      "@       @              @      "@      @      @              @      @               @      @      @      �?       @      �?                       @      @      �?      �?              @      �?       @              �?      �?              �?      �?              �?             Pq@     �C@     �p@     �B@     �j@      A@     �f@      ?@      "@      @       @      @       @      @      �?      @      �?      @      �?                      @              �?      �?                      @      @             �e@      8@     @X@      @     @T@      @      1@              P@      @      <@       @       @      �?              �?       @              :@      �?      *@              *@      �?      @              $@      �?      "@      �?      �?              B@      �?      &@              9@      �?      "@      �?       @              �?      �?      0@              0@      @              �?      0@       @      @      �?              �?      @              (@      �?      @      �?      @                      �?       @             �R@      2@     �R@      0@      7@      �?      $@              *@      �?      @      �?      @              �?      �?              �?      �?              "@              J@      .@      @      �?              �?      @              G@      ,@      2@      @      "@      @      @      @       @       @       @      �?      @              "@              <@      &@               @      <@      "@      .@              *@      "@      @      "@              @      @      @               @      @       @      @      �?      @              �?      �?              �?      @                       @     �@@      @       @              9@      @      @       @      @      �?      @               @      �?              �?       @                      �?      2@      �?      ,@              @      �?       @               @      �?              �?       @             �K@      @     �I@       @      I@       @      4@              >@       @      @              ;@       @      @       @      @      �?      @                      �?      @      �?      @                      �?      4@              �?              @      �?      �?      �?              �?      �?              @               @       @      @              @       @      �?       @      �?                       @      @                       @      L@      8@     �J@      8@       @      *@       @      $@              $@       @                      @     �F@      &@      @@      &@      �?      @      �?      �?              �?      �?                      @      ?@      @      (@              3@      @      @      @               @      @      @      @       @      @              @       @               @      @                       @      *@              *@              @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�%hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM1huh*h-K ��h/��R�(KM1��h|�B@L                             @
Ϛ����?�           @�@                                  �C@���!pc�?             F@                                   @��G���?            �B@        ������������������������       �                     *@               
                    @�q�q�?             8@              	                    �?��S�ۿ?             .@                               P��%@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     @                                ��T?@�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @                                   @����X�?             @       ������������������������       �                     @        ������������������������       �                      @               N                    �?�'���?�           ��@               !                 ��K.@�`���?C            �X@                                   P,@������?            �B@                                   @PN��T'�?             ;@        ������������������������       �                     �?                                  @@ȵHPS!�?             :@                                  �?�S����?             3@        ������������������������       �                     �?                                ���@�����H�?             2@        ������������������������       �                     @                                   �?8�Z$���?             *@                                  5@z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@        "       K                 �\@�jTM��?,            �N@       #       ,                    �?f.i��n�?$            �F@        $       +                     �?P���Q�?             4@       %       *                    �?$�q-�?             *@       &       '                   �G@ףp=
�?             $@       ������������������������       �                      @        (       )                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        -       <                    �?�q�����?             9@       .       ;                    �?��S���?             .@       /       :                  �}S@�q�q�?
             (@       0       9                      @���|���?	             &@       1       2                   �;@���Q��?             $@        ������������������������       �                      @        3       4                 �ܵ<@      �?              @        ������������������������       �                      @        5       8                   �B@�q�q�?             @       6       7                   �L@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        =       F                   �C@      �?	             $@       >       E                   �:@�q�q�?             @       ?       @                 H�<@      �?             @        ������������������������       �                     �?        A       D                     �?�q�q�?             @       B       C                 8�T@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        G       H                   @H@      �?             @        ������������������������       �                     �?        I       J                 ���X@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        L       M                   �6@      �?             0@        ������������������������       �                     �?        ������������������������       �                     .@        O                        x#J@��h!��?l           Ё@       P       �                 `f�$@�l�6���?6           �~@       Q       �                    @P��S�I�?�             q@       R       m                    �?(5DSbq�?�             q@        S       l                    �?8�A�0��?             F@       T       k                    �?��
ц��?            �C@       U       j                 pF @��+��?            �B@       V       _                    �?�q�q�?             ;@       W       X                   �2@d}h���?
             ,@        ������������������������       �                     @        Y       ^                 �&B@���!pc�?             &@       Z       [                   �8@      �?              @        ������������������������       �                     �?        \       ]                 ���@����X�?             @        ������������������������       �                      @        ������������������������       ����Q��?             @        ������������������������       �                     @        `       i                   �9@��
ц��?	             *@       a       h                   �6@�q�q�?             "@       b       c                 ���@���Q��?             @        ������������������������       �                      @        d       g                 �&B@�q�q�?             @       e       f                    4@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                      @        ������������������������       �                     @        n       y                 ��@@݈g>h�?�            �l@        o       t                   �8@ 7���B�?/            @T@        p       s                 ���@�KM�]�?             3@        q       r                    7@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     *@        u       v                  ��@0�z��?�?#             O@       ������������������������       �                    �G@        w       x                    >@��S�ۿ?
             .@       ������������������������       �ףp=
�?             $@        ������������������������       �                     @        z       �                    �?�q��/��?Z            `b@       {       �                   @@@(N:!���?U            �a@       |       �                   �:@؇���X�??            @Z@        }       �                   �3@HP�s��?             I@        ~       �                   �2@�J�4�?             9@              �                 ��Y @�C��2(�?	             &@        �       �                 pf�@z�G�z�?             @        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     @        �       �                 �?�@d}h���?             ,@        ������������������������       �                     @        �       �                 `�8"@և���X�?             @       ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     9@        �       �                 pb@z�G�z�?!            �K@        �       �                   �=@և���X�?             @       �       �                   �;@�q�q�?             @        ������������������������       �                     �?        �       �                 �?$@���Q��?             @       ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �;@8��8���?             H@        ������������������������       �                     �?        �       �                 ��) @��E�B��?            �G@       �       �                 �?�@      �?             @@       ������������������������       �                     .@        �       �                    ?@�t����?             1@       ������������������������       �                     .@        ������������������������       �                      @        �       �                 ��y @������?             .@        ������������������������       �                      @        �       �                   �>@8�Z$���?             *@       �       �                   �<@      �?              @       ������������������������       �                     @        �       �                 ���"@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                   @C@��?^�k�?            �A@        ������������������������       �                     4@        �       �                   �C@��S�ۿ?             .@        ������������������������       ��q�q�?             @        ������������������������       �        	             (@        �       �                    �?����X�?             @       �       �                    �?���Q��?             @        �       �                   �9@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?�h^���?�            �k@        �       �                    @H�z���?7             T@       �       �                    �?x!'ǯ�?3            �R@       �       �                    �?�:�B��?*            �M@        ������������������������       �                     @        �       �                   �?@r�����?&            �J@       �       �                     @�q�q�?             ;@       �       �                    6@r�q��?             2@        �       �                   �;@�z�G��?             $@       �       �                    �?      �?             @       �       �                   �6@���Q��?             @        ������������������������       �                     �?        ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�q�q�?             "@        �       �                 ��1@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �? ��WV�?             :@       ������������������������       �                     3@        �       �                 `f�/@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ���B@�q�q�?	             .@       �       �                    @�θ�?             *@       �       �                 0339@�z�G��?             $@       �       �                 @34@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �                          �?�{"z;m�?X            �a@       �                           �? �Cc}�?E             \@       �       �                   �R@d/
k�?C             [@       �       �                    �?��hq��?B            �Z@       �       �                    �?��Lɿ��?4            �T@        ������������������������       �                      @        �       �                     �?�����H�?2            @T@        �       �                   �>@�+e�X�?             9@       �       �                   �J@��
ц��?
             *@       �       �                 `fF:@      �?              @        ������������������������       �                     �?        �       �                 `f�;@؇���X�?             @        ������������������������       �                     @        �       �                   `B@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        �       �                    4@�h����?              L@        �       �                    &@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �*@@9G��?            �H@       �       �                   �@@ >�֕�?            �A@        ������������������������       �                     1@        �       �                   @A@�����H�?             2@        ������������������������       �      �?              @        �       �                 `f�)@      �?	             0@        ������������������������       �                      @        �       �                   @D@      �?              @        ������������������������       �                     @        �       �                   �F@z�G�z�?             @        ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �        	             ,@        �       �                   �?@ �q�q�?             8@        ������������������������       �                     (@        �       �                   �:@�8��8��?             (@       �       �                   �7@�����H�?             "@        ������������������������       �                      @        �       �                    C@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?                                 �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @                                 0@XB���?             =@                                 �?؇���X�?             @        ������������������������       �                     @                                 �?      �?             @        ������������������������       �                     �?        	      
                  �5@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     6@                                 �?L�qA��?6            �R@                                �?��-�=��?            �C@        ������������������������       �                      @                                 @������?            �B@                               �:@ >�֕�?            �A@                              ���`@؇���X�?	             ,@       ������������������������       �                     "@                                �8@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     5@        ������������������������       �                      @              ,                   �?�q�q�?             B@                                �?�\��N��?             3@                                 >@؇���X�?             @                                ;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                     @               !                   7@      �?	             (@        ������������������������       �                      @        "      )                   �?�z�G��?             $@       #      $                   <@      �?              @        ������������������������       �                     �?        %      (                  �D@؇���X�?             @       &      '                03U@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        *      +                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        -      0                  @F@@�0�!��?
             1@       .      /                   @@�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �t�bh�h*h-K ��h/��R�(KM1KK��h]�B       `}@     @n@      (@      @@      @      >@              *@      @      1@      �?      ,@      �?      "@      �?                      "@              @      @      @      @                      @      @       @      @                       @     �|@     @j@      H@      I@     �@@      @      7@      @              �?      7@      @      0@      @              �?      0@       @      @              &@       @       @       @               @       @              @              @              $@              .@      G@      ,@      ?@      �?      3@      �?      (@      �?      "@               @      �?      �?      �?                      �?              @              @      *@      (@       @      @      @      @      @      @      @      @               @      @      @       @               @      @      �?      @              @      �?              �?                      �?      �?              @              @      @      @       @       @       @              �?       @      �?      �?      �?              �?      �?              �?               @              �?      @              �?      �?       @               @      �?              �?      .@      �?                      .@     �y@      d@     �w@     @\@      m@     �D@      m@     �C@      :@      2@      5@      2@      3@      2@      "@      2@      @      &@              @      @       @      @      @      �?               @      @               @       @      @              @      @      @      @      @       @      @               @       @      �?      �?      �?      �?                      �?      �?              @                      @      $@               @              @             �i@      5@     �S@      @      1@       @      @       @      @                       @      *@             �N@      �?     �G@              ,@      �?      "@      �?      @              `@      2@      _@      0@     �V@      .@      G@      @      5@      @      $@      �?      @      �?      @              �?      �?      @              &@      @      @              @      @      �?      @      @              9@              F@      &@      @      @       @      @              �?       @      @      �?      @      �?              �?             �D@      @              �?     �D@      @      >@       @      .@              .@       @      .@                       @      &@      @               @      &@       @      @       @      @               @       @       @                       @      @              A@      �?      4@              ,@      �?       @      �?      (@              @       @      @       @      �?       @               @      �?               @               @                       @     �b@      R@      5@     �M@      .@     �M@      $@     �H@              @      $@     �E@      "@      2@      @      .@      @      @      @      @       @      @              �?       @       @      �?                      @               @      @      @       @      @              @       @              @              �?      9@              3@      �?      @      �?                      @      @      $@      @      $@      @      @      @       @               @      @                      @              @       @              @              `@      *@      Y@      (@     @X@      &@     @X@      $@     �R@      "@       @              R@      "@      3@      @      @      @       @      @      �?              �?      @              @      �?       @               @      �?              @              (@             �J@      @      @      �?              �?      @             �G@       @     �@@       @      1@              0@       @      �?      �?      .@      �?       @              @      �?      @              @      �?       @      �?       @              ,@              7@      �?      (@              &@      �?       @      �?       @              @      �?              �?      @              @                      �?      @      �?              �?      @              <@      �?      @      �?      @              @      �?      �?               @      �?              �?       @              6@              <@     �G@      @     �A@               @      @     �@@       @     �@@       @      (@              "@       @      @              @       @                      5@       @              8@      (@      $@      "@      �?      @      �?       @              �?      �?      �?              @      "@      @       @              @      @      @       @              �?      @      �?       @      �?       @                      �?      @              �?      �?      �?                      �?      ,@      @      @      @      @                      @       @        �t�bubhhubehhub.